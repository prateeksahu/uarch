module test_all;

	reg	[7:0]	inst_bytes	[781:0][11:0];
	reg	[3:0]	inst_size	[781:0];

	initial 
	begin

		inst_bytes	[0][0]	= 8'h04;
		inst_bytes	[0][1]	= 8'h11;
		inst_size	[0]		= 4'd2;

		inst_bytes	[1][0]	= 8'h66;
		inst_bytes	[1][1]	= 8'h05;
		inst_bytes	[1][2]	= 8'h11;
		inst_bytes	[1][3]	= 8'h12;
		inst_size	[1]		= 4'd4;

		inst_bytes	[2][0]	= 8'h05;
		inst_bytes	[2][1]	= 8'h11;
		inst_bytes	[2][2]	= 8'h12;
		inst_bytes	[2][3]	= 8'h13;
		inst_bytes	[2][4]	= 8'h14;
		inst_size	[2]		= 4'd5;

		inst_bytes	[3][0]	= 8'h80;
		inst_bytes	[3][1]	= 8'h01;
		inst_bytes	[3][2]	= 8'h11;
		inst_size	[3]		= 4'd3;

		inst_bytes	[4][0]	= 8'h80;
		inst_bytes	[4][1]	= 8'h04;
		inst_bytes	[4][2]	= 8'h52;
		inst_bytes	[4][3]	= 8'h11;
		inst_size	[4]		= 4'd4;

		inst_bytes	[5][0]	= 8'h80;
		inst_bytes	[5][1]	= 8'h05;
		inst_bytes	[5][2]	= 8'h01;
		inst_bytes	[5][3]	= 8'h02;
		inst_bytes	[5][4]	= 8'h03;
		inst_bytes	[5][5]	= 8'h04;
		inst_bytes	[5][6]	= 8'h11;
		inst_size	[5]		= 4'd7;

		inst_bytes	[6][0]	= 8'h80;
		inst_bytes	[6][1]	= 8'h41;
		inst_bytes	[6][2]	= 8'h01;
		inst_bytes	[6][3]	= 8'h11;
		inst_size	[6]		= 4'd4;

		inst_bytes	[7][0]	= 8'h80;
		inst_bytes	[7][1]	= 8'h44;
		inst_bytes	[7][2]	= 8'h52;
		inst_bytes	[7][3]	= 8'h01;
		inst_bytes	[7][4]	= 8'h11;
		inst_size	[7]		= 4'd5;

		inst_bytes	[8][0]	= 8'h80;
		inst_bytes	[8][1]	= 8'h81;
		inst_bytes	[8][2]	= 8'h01;
		inst_bytes	[8][3]	= 8'h02;
		inst_bytes	[8][4]	= 8'h03;
		inst_bytes	[8][5]	= 8'h04;
		inst_bytes	[8][6]	= 8'h11;
		inst_size	[8]		= 4'd7;

		inst_bytes	[9][0]	= 8'h80;
		inst_bytes	[9][1]	= 8'h84;
		inst_bytes	[9][2]	= 8'h52;
		inst_bytes	[9][3]	= 8'h01;
		inst_bytes	[9][4]	= 8'h02;
		inst_bytes	[9][5]	= 8'h03;
		inst_bytes	[9][6]	= 8'h04;
		inst_bytes	[9][7]	= 8'h11;
		inst_size	[9]		= 4'd8;

		inst_bytes	[10][0]	= 8'h80;
		inst_bytes	[10][1]	= 8'hC1;
		inst_bytes	[10][2]	= 8'h11;
		inst_size	[10]		= 4'd3;

		inst_bytes	[11][0]	= 8'h66;
		inst_bytes	[11][1]	= 8'h81;
		inst_bytes	[11][2]	= 8'h01;
		inst_bytes	[11][3]	= 8'h11;
		inst_bytes	[11][4]	= 8'h12;
		inst_size	[11]		= 4'd5;

		inst_bytes	[12][0]	= 8'h66;
		inst_bytes	[12][1]	= 8'h81;
		inst_bytes	[12][2]	= 8'h04;
		inst_bytes	[12][3]	= 8'h52;
		inst_bytes	[12][4]	= 8'h11;
		inst_bytes	[12][5]	= 8'h12;
		inst_size	[12]		= 4'd6;

		inst_bytes	[13][0]	= 8'h66;
		inst_bytes	[13][1]	= 8'h81;
		inst_bytes	[13][2]	= 8'h05;
		inst_bytes	[13][3]	= 8'h01;
		inst_bytes	[13][4]	= 8'h02;
		inst_bytes	[13][5]	= 8'h03;
		inst_bytes	[13][6]	= 8'h04;
		inst_bytes	[13][7]	= 8'h11;
		inst_bytes	[13][8]	= 8'h12;
		inst_size	[13]		= 4'd9;

		inst_bytes	[14][0]	= 8'h66;
		inst_bytes	[14][1]	= 8'h81;
		inst_bytes	[14][2]	= 8'h41;
		inst_bytes	[14][3]	= 8'h01;
		inst_bytes	[14][4]	= 8'h11;
		inst_bytes	[14][5]	= 8'h12;
		inst_size	[14]		= 4'd6;

		inst_bytes	[15][0]	= 8'h66;
		inst_bytes	[15][1]	= 8'h81;
		inst_bytes	[15][2]	= 8'h44;
		inst_bytes	[15][3]	= 8'h52;
		inst_bytes	[15][4]	= 8'h01;
		inst_bytes	[15][5]	= 8'h11;
		inst_bytes	[15][6]	= 8'h12;
		inst_size	[15]		= 4'd7;

		inst_bytes	[16][0]	= 8'h66;
		inst_bytes	[16][1]	= 8'h81;
		inst_bytes	[16][2]	= 8'h81;
		inst_bytes	[16][3]	= 8'h01;
		inst_bytes	[16][4]	= 8'h02;
		inst_bytes	[16][5]	= 8'h03;
		inst_bytes	[16][6]	= 8'h04;
		inst_bytes	[16][7]	= 8'h11;
		inst_bytes	[16][8]	= 8'h12;
		inst_size	[16]		= 4'd9;

		inst_bytes	[17][0]	= 8'h66;
		inst_bytes	[17][1]	= 8'h81;
		inst_bytes	[17][2]	= 8'h84;
		inst_bytes	[17][3]	= 8'h52;
		inst_bytes	[17][4]	= 8'h01;
		inst_bytes	[17][5]	= 8'h02;
		inst_bytes	[17][6]	= 8'h03;
		inst_bytes	[17][7]	= 8'h04;
		inst_bytes	[17][8]	= 8'h11;
		inst_bytes	[17][9]	= 8'h12;
		inst_size	[17]		= 4'd10;

		inst_bytes	[18][0]	= 8'h66;
		inst_bytes	[18][1]	= 8'h81;
		inst_bytes	[18][2]	= 8'hC1;
		inst_bytes	[18][3]	= 8'h11;
		inst_bytes	[18][4]	= 8'h12;
		inst_size	[18]		= 4'd5;

		inst_bytes	[19][0]	= 8'h81;
		inst_bytes	[19][1]	= 8'h01;
		inst_bytes	[19][2]	= 8'h11;
		inst_bytes	[19][3]	= 8'h12;
		inst_bytes	[19][4]	= 8'h13;
		inst_bytes	[19][5]	= 8'h14;
		inst_size	[19]		= 4'd6;

		inst_bytes	[20][0]	= 8'h81;
		inst_bytes	[20][1]	= 8'h04;
		inst_bytes	[20][2]	= 8'h52;
		inst_bytes	[20][3]	= 8'h11;
		inst_bytes	[20][4]	= 8'h12;
		inst_bytes	[20][5]	= 8'h13;
		inst_bytes	[20][6]	= 8'h14;
		inst_size	[20]		= 4'd7;

		inst_bytes	[21][0]	= 8'h81;
		inst_bytes	[21][1]	= 8'h05;
		inst_bytes	[21][2]	= 8'h01;
		inst_bytes	[21][3]	= 8'h02;
		inst_bytes	[21][4]	= 8'h03;
		inst_bytes	[21][5]	= 8'h04;
		inst_bytes	[21][6]	= 8'h11;
		inst_bytes	[21][7]	= 8'h12;
		inst_bytes	[21][8]	= 8'h13;
		inst_bytes	[21][9]	= 8'h14;
		inst_size	[21]		= 4'd10;

		inst_bytes	[22][0]	= 8'h81;
		inst_bytes	[22][1]	= 8'h41;
		inst_bytes	[22][2]	= 8'h01;
		inst_bytes	[22][3]	= 8'h11;
		inst_bytes	[22][4]	= 8'h12;
		inst_bytes	[22][5]	= 8'h13;
		inst_bytes	[22][6]	= 8'h14;
		inst_size	[22]		= 4'd7;

		inst_bytes	[23][0]	= 8'h81;
		inst_bytes	[23][1]	= 8'h44;
		inst_bytes	[23][2]	= 8'h52;
		inst_bytes	[23][3]	= 8'h01;
		inst_bytes	[23][4]	= 8'h11;
		inst_bytes	[23][5]	= 8'h12;
		inst_bytes	[23][6]	= 8'h13;
		inst_bytes	[23][7]	= 8'h14;
		inst_size	[23]		= 4'd8;

		inst_bytes	[24][0]	= 8'h81;
		inst_bytes	[24][1]	= 8'h81;
		inst_bytes	[24][2]	= 8'h01;
		inst_bytes	[24][3]	= 8'h02;
		inst_bytes	[24][4]	= 8'h03;
		inst_bytes	[24][5]	= 8'h04;
		inst_bytes	[24][6]	= 8'h11;
		inst_bytes	[24][7]	= 8'h12;
		inst_bytes	[24][8]	= 8'h13;
		inst_bytes	[24][9]	= 8'h14;
		inst_size	[24]		= 4'd10;

		inst_bytes	[25][0]	= 8'h81;
		inst_bytes	[25][1]	= 8'h84;
		inst_bytes	[25][2]	= 8'h52;
		inst_bytes	[25][3]	= 8'h01;
		inst_bytes	[25][4]	= 8'h02;
		inst_bytes	[25][5]	= 8'h03;
		inst_bytes	[25][6]	= 8'h04;
		inst_bytes	[25][7]	= 8'h11;
		inst_bytes	[25][8]	= 8'h12;
		inst_bytes	[25][9]	= 8'h13;
		inst_bytes	[25][10]	= 8'h14;
		inst_size	[25]		= 4'd11;

		inst_bytes	[26][0]	= 8'h81;
		inst_bytes	[26][1]	= 8'hC1;
		inst_bytes	[26][2]	= 8'h11;
		inst_bytes	[26][3]	= 8'h12;
		inst_bytes	[26][4]	= 8'h13;
		inst_bytes	[26][5]	= 8'h14;
		inst_size	[26]		= 4'd6;

		inst_bytes	[27][0]	= 8'h83;
		inst_bytes	[27][1]	= 8'h01;
		inst_bytes	[27][2]	= 8'h11;
		inst_size	[27]		= 4'd3;

		inst_bytes	[28][0]	= 8'h83;
		inst_bytes	[28][1]	= 8'h04;
		inst_bytes	[28][2]	= 8'h52;
		inst_bytes	[28][3]	= 8'h11;
		inst_size	[28]		= 4'd4;

		inst_bytes	[29][0]	= 8'h83;
		inst_bytes	[29][1]	= 8'h05;
		inst_bytes	[29][2]	= 8'h01;
		inst_bytes	[29][3]	= 8'h02;
		inst_bytes	[29][4]	= 8'h03;
		inst_bytes	[29][5]	= 8'h04;
		inst_bytes	[29][6]	= 8'h11;
		inst_size	[29]		= 4'd7;

		inst_bytes	[30][0]	= 8'h83;
		inst_bytes	[30][1]	= 8'h41;
		inst_bytes	[30][2]	= 8'h01;
		inst_bytes	[30][3]	= 8'h11;
		inst_size	[30]		= 4'd4;

		inst_bytes	[31][0]	= 8'h83;
		inst_bytes	[31][1]	= 8'h44;
		inst_bytes	[31][2]	= 8'h52;
		inst_bytes	[31][3]	= 8'h01;
		inst_bytes	[31][4]	= 8'h11;
		inst_size	[31]		= 4'd5;

		inst_bytes	[32][0]	= 8'h83;
		inst_bytes	[32][1]	= 8'h81;
		inst_bytes	[32][2]	= 8'h01;
		inst_bytes	[32][3]	= 8'h02;
		inst_bytes	[32][4]	= 8'h03;
		inst_bytes	[32][5]	= 8'h04;
		inst_bytes	[32][6]	= 8'h11;
		inst_size	[32]		= 4'd7;

		inst_bytes	[33][0]	= 8'h83;
		inst_bytes	[33][1]	= 8'h84;
		inst_bytes	[33][2]	= 8'h52;
		inst_bytes	[33][3]	= 8'h01;
		inst_bytes	[33][4]	= 8'h02;
		inst_bytes	[33][5]	= 8'h03;
		inst_bytes	[33][6]	= 8'h04;
		inst_bytes	[33][7]	= 8'h11;
		inst_size	[33]		= 4'd8;

		inst_bytes	[34][0]	= 8'h83;
		inst_bytes	[34][1]	= 8'hC1;
		inst_bytes	[34][2]	= 8'h11;
		inst_size	[34]		= 4'd3;

		inst_bytes	[35][0]	= 8'h83;
		inst_bytes	[35][1]	= 8'h01;
		inst_bytes	[35][2]	= 8'h11;
		inst_size	[35]		= 4'd3;

		inst_bytes	[36][0]	= 8'h83;
		inst_bytes	[36][1]	= 8'h04;
		inst_bytes	[36][2]	= 8'h52;
		inst_bytes	[36][3]	= 8'h11;
		inst_size	[36]		= 4'd4;

		inst_bytes	[37][0]	= 8'h83;
		inst_bytes	[37][1]	= 8'h05;
		inst_bytes	[37][2]	= 8'h01;
		inst_bytes	[37][3]	= 8'h02;
		inst_bytes	[37][4]	= 8'h03;
		inst_bytes	[37][5]	= 8'h04;
		inst_bytes	[37][6]	= 8'h11;
		inst_size	[37]		= 4'd7;

		inst_bytes	[38][0]	= 8'h83;
		inst_bytes	[38][1]	= 8'h41;
		inst_bytes	[38][2]	= 8'h01;
		inst_bytes	[38][3]	= 8'h11;
		inst_size	[38]		= 4'd4;

		inst_bytes	[39][0]	= 8'h83;
		inst_bytes	[39][1]	= 8'h44;
		inst_bytes	[39][2]	= 8'h52;
		inst_bytes	[39][3]	= 8'h01;
		inst_bytes	[39][4]	= 8'h11;
		inst_size	[39]		= 4'd5;

		inst_bytes	[40][0]	= 8'h83;
		inst_bytes	[40][1]	= 8'h81;
		inst_bytes	[40][2]	= 8'h01;
		inst_bytes	[40][3]	= 8'h02;
		inst_bytes	[40][4]	= 8'h03;
		inst_bytes	[40][5]	= 8'h04;
		inst_bytes	[40][6]	= 8'h11;
		inst_size	[40]		= 4'd7;

		inst_bytes	[41][0]	= 8'h83;
		inst_bytes	[41][1]	= 8'h84;
		inst_bytes	[41][2]	= 8'h52;
		inst_bytes	[41][3]	= 8'h01;
		inst_bytes	[41][4]	= 8'h02;
		inst_bytes	[41][5]	= 8'h03;
		inst_bytes	[41][6]	= 8'h04;
		inst_bytes	[41][7]	= 8'h11;
		inst_size	[41]		= 4'd8;

		inst_bytes	[42][0]	= 8'h83;
		inst_bytes	[42][1]	= 8'hC1;
		inst_bytes	[42][2]	= 8'h11;
		inst_size	[42]		= 4'd3;

		inst_bytes	[43][0]	= 8'h00;
		inst_bytes	[43][1]	= 8'h01;
		inst_size	[43]		= 4'd2;

		inst_bytes	[44][0]	= 8'h00;
		inst_bytes	[44][1]	= 8'h04;
		inst_bytes	[44][2]	= 8'h52;
		inst_size	[44]		= 4'd3;

		inst_bytes	[45][0]	= 8'h00;
		inst_bytes	[45][1]	= 8'h05;
		inst_bytes	[45][2]	= 8'h01;
		inst_bytes	[45][3]	= 8'h02;
		inst_bytes	[45][4]	= 8'h03;
		inst_bytes	[45][5]	= 8'h04;
		inst_size	[45]		= 4'd6;

		inst_bytes	[46][0]	= 8'h00;
		inst_bytes	[46][1]	= 8'h41;
		inst_bytes	[46][2]	= 8'h01;
		inst_size	[46]		= 4'd3;

		inst_bytes	[47][0]	= 8'h00;
		inst_bytes	[47][1]	= 8'h44;
		inst_bytes	[47][2]	= 8'h52;
		inst_bytes	[47][3]	= 8'h01;
		inst_size	[47]		= 4'd4;

		inst_bytes	[48][0]	= 8'h00;
		inst_bytes	[48][1]	= 8'h81;
		inst_bytes	[48][2]	= 8'h01;
		inst_bytes	[48][3]	= 8'h02;
		inst_bytes	[48][4]	= 8'h03;
		inst_bytes	[48][5]	= 8'h04;
		inst_size	[48]		= 4'd6;

		inst_bytes	[49][0]	= 8'h00;
		inst_bytes	[49][1]	= 8'h84;
		inst_bytes	[49][2]	= 8'h52;
		inst_bytes	[49][3]	= 8'h01;
		inst_bytes	[49][4]	= 8'h02;
		inst_bytes	[49][5]	= 8'h03;
		inst_bytes	[49][6]	= 8'h04;
		inst_size	[49]		= 4'd7;

		inst_bytes	[50][0]	= 8'h00;
		inst_bytes	[50][1]	= 8'hC1;
		inst_size	[50]		= 4'd2;

		inst_bytes	[51][0]	= 8'h01;
		inst_bytes	[51][1]	= 8'h01;
		inst_size	[51]		= 4'd2;

		inst_bytes	[52][0]	= 8'h01;
		inst_bytes	[52][1]	= 8'h04;
		inst_bytes	[52][2]	= 8'h52;
		inst_size	[52]		= 4'd3;

		inst_bytes	[53][0]	= 8'h01;
		inst_bytes	[53][1]	= 8'h05;
		inst_bytes	[53][2]	= 8'h01;
		inst_bytes	[53][3]	= 8'h02;
		inst_bytes	[53][4]	= 8'h03;
		inst_bytes	[53][5]	= 8'h04;
		inst_size	[53]		= 4'd6;

		inst_bytes	[54][0]	= 8'h01;
		inst_bytes	[54][1]	= 8'h41;
		inst_bytes	[54][2]	= 8'h01;
		inst_size	[54]		= 4'd3;

		inst_bytes	[55][0]	= 8'h01;
		inst_bytes	[55][1]	= 8'h44;
		inst_bytes	[55][2]	= 8'h52;
		inst_bytes	[55][3]	= 8'h01;
		inst_size	[55]		= 4'd4;

		inst_bytes	[56][0]	= 8'h01;
		inst_bytes	[56][1]	= 8'h81;
		inst_bytes	[56][2]	= 8'h01;
		inst_bytes	[56][3]	= 8'h02;
		inst_bytes	[56][4]	= 8'h03;
		inst_bytes	[56][5]	= 8'h04;
		inst_size	[56]		= 4'd6;

		inst_bytes	[57][0]	= 8'h01;
		inst_bytes	[57][1]	= 8'h84;
		inst_bytes	[57][2]	= 8'h52;
		inst_bytes	[57][3]	= 8'h01;
		inst_bytes	[57][4]	= 8'h02;
		inst_bytes	[57][5]	= 8'h03;
		inst_bytes	[57][6]	= 8'h04;
		inst_size	[57]		= 4'd7;

		inst_bytes	[58][0]	= 8'h01;
		inst_bytes	[58][1]	= 8'hC1;
		inst_size	[58]		= 4'd2;

		inst_bytes	[59][0]	= 8'h01;
		inst_bytes	[59][1]	= 8'h01;
		inst_size	[59]		= 4'd2;

		inst_bytes	[60][0]	= 8'h01;
		inst_bytes	[60][1]	= 8'h04;
		inst_bytes	[60][2]	= 8'h52;
		inst_size	[60]		= 4'd3;

		inst_bytes	[61][0]	= 8'h01;
		inst_bytes	[61][1]	= 8'h05;
		inst_bytes	[61][2]	= 8'h01;
		inst_bytes	[61][3]	= 8'h02;
		inst_bytes	[61][4]	= 8'h03;
		inst_bytes	[61][5]	= 8'h04;
		inst_size	[61]		= 4'd6;

		inst_bytes	[62][0]	= 8'h01;
		inst_bytes	[62][1]	= 8'h41;
		inst_bytes	[62][2]	= 8'h01;
		inst_size	[62]		= 4'd3;

		inst_bytes	[63][0]	= 8'h01;
		inst_bytes	[63][1]	= 8'h44;
		inst_bytes	[63][2]	= 8'h52;
		inst_bytes	[63][3]	= 8'h01;
		inst_size	[63]		= 4'd4;

		inst_bytes	[64][0]	= 8'h01;
		inst_bytes	[64][1]	= 8'h81;
		inst_bytes	[64][2]	= 8'h01;
		inst_bytes	[64][3]	= 8'h02;
		inst_bytes	[64][4]	= 8'h03;
		inst_bytes	[64][5]	= 8'h04;
		inst_size	[64]		= 4'd6;

		inst_bytes	[65][0]	= 8'h01;
		inst_bytes	[65][1]	= 8'h84;
		inst_bytes	[65][2]	= 8'h52;
		inst_bytes	[65][3]	= 8'h01;
		inst_bytes	[65][4]	= 8'h02;
		inst_bytes	[65][5]	= 8'h03;
		inst_bytes	[65][6]	= 8'h04;
		inst_size	[65]		= 4'd7;

		inst_bytes	[66][0]	= 8'h01;
		inst_bytes	[66][1]	= 8'hC1;
		inst_size	[66]		= 4'd2;

		inst_bytes	[67][0]	= 8'h02;
		inst_bytes	[67][1]	= 8'h01;
		inst_size	[67]		= 4'd2;

		inst_bytes	[68][0]	= 8'h02;
		inst_bytes	[68][1]	= 8'h04;
		inst_bytes	[68][2]	= 8'h52;
		inst_size	[68]		= 4'd3;

		inst_bytes	[69][0]	= 8'h02;
		inst_bytes	[69][1]	= 8'h05;
		inst_bytes	[69][2]	= 8'h01;
		inst_bytes	[69][3]	= 8'h02;
		inst_bytes	[69][4]	= 8'h03;
		inst_bytes	[69][5]	= 8'h04;
		inst_size	[69]		= 4'd6;

		inst_bytes	[70][0]	= 8'h02;
		inst_bytes	[70][1]	= 8'h41;
		inst_bytes	[70][2]	= 8'h01;
		inst_size	[70]		= 4'd3;

		inst_bytes	[71][0]	= 8'h02;
		inst_bytes	[71][1]	= 8'h44;
		inst_bytes	[71][2]	= 8'h52;
		inst_bytes	[71][3]	= 8'h01;
		inst_size	[71]		= 4'd4;

		inst_bytes	[72][0]	= 8'h02;
		inst_bytes	[72][1]	= 8'h81;
		inst_bytes	[72][2]	= 8'h01;
		inst_bytes	[72][3]	= 8'h02;
		inst_bytes	[72][4]	= 8'h03;
		inst_bytes	[72][5]	= 8'h04;
		inst_size	[72]		= 4'd6;

		inst_bytes	[73][0]	= 8'h02;
		inst_bytes	[73][1]	= 8'h84;
		inst_bytes	[73][2]	= 8'h52;
		inst_bytes	[73][3]	= 8'h01;
		inst_bytes	[73][4]	= 8'h02;
		inst_bytes	[73][5]	= 8'h03;
		inst_bytes	[73][6]	= 8'h04;
		inst_size	[73]		= 4'd7;

		inst_bytes	[74][0]	= 8'h02;
		inst_bytes	[74][1]	= 8'hC1;
		inst_size	[74]		= 4'd2;

		inst_bytes	[75][0]	= 8'h03;
		inst_bytes	[75][1]	= 8'h01;
		inst_size	[75]		= 4'd2;

		inst_bytes	[76][0]	= 8'h03;
		inst_bytes	[76][1]	= 8'h04;
		inst_bytes	[76][2]	= 8'h52;
		inst_size	[76]		= 4'd3;

		inst_bytes	[77][0]	= 8'h03;
		inst_bytes	[77][1]	= 8'h05;
		inst_bytes	[77][2]	= 8'h01;
		inst_bytes	[77][3]	= 8'h02;
		inst_bytes	[77][4]	= 8'h03;
		inst_bytes	[77][5]	= 8'h04;
		inst_size	[77]		= 4'd6;

		inst_bytes	[78][0]	= 8'h03;
		inst_bytes	[78][1]	= 8'h41;
		inst_bytes	[78][2]	= 8'h01;
		inst_size	[78]		= 4'd3;

		inst_bytes	[79][0]	= 8'h03;
		inst_bytes	[79][1]	= 8'h44;
		inst_bytes	[79][2]	= 8'h52;
		inst_bytes	[79][3]	= 8'h01;
		inst_size	[79]		= 4'd4;

		inst_bytes	[80][0]	= 8'h03;
		inst_bytes	[80][1]	= 8'h81;
		inst_bytes	[80][2]	= 8'h01;
		inst_bytes	[80][3]	= 8'h02;
		inst_bytes	[80][4]	= 8'h03;
		inst_bytes	[80][5]	= 8'h04;
		inst_size	[80]		= 4'd6;

		inst_bytes	[81][0]	= 8'h03;
		inst_bytes	[81][1]	= 8'h84;
		inst_bytes	[81][2]	= 8'h52;
		inst_bytes	[81][3]	= 8'h01;
		inst_bytes	[81][4]	= 8'h02;
		inst_bytes	[81][5]	= 8'h03;
		inst_bytes	[81][6]	= 8'h04;
		inst_size	[81]		= 4'd7;

		inst_bytes	[82][0]	= 8'h03;
		inst_bytes	[82][1]	= 8'hC1;
		inst_size	[82]		= 4'd2;

		inst_bytes	[83][0]	= 8'h03;
		inst_bytes	[83][1]	= 8'h01;
		inst_size	[83]		= 4'd2;

		inst_bytes	[84][0]	= 8'h03;
		inst_bytes	[84][1]	= 8'h04;
		inst_bytes	[84][2]	= 8'h52;
		inst_size	[84]		= 4'd3;

		inst_bytes	[85][0]	= 8'h03;
		inst_bytes	[85][1]	= 8'h05;
		inst_bytes	[85][2]	= 8'h01;
		inst_bytes	[85][3]	= 8'h02;
		inst_bytes	[85][4]	= 8'h03;
		inst_bytes	[85][5]	= 8'h04;
		inst_size	[85]		= 4'd6;

		inst_bytes	[86][0]	= 8'h03;
		inst_bytes	[86][1]	= 8'h41;
		inst_bytes	[86][2]	= 8'h01;
		inst_size	[86]		= 4'd3;

		inst_bytes	[87][0]	= 8'h03;
		inst_bytes	[87][1]	= 8'h44;
		inst_bytes	[87][2]	= 8'h52;
		inst_bytes	[87][3]	= 8'h01;
		inst_size	[87]		= 4'd4;

		inst_bytes	[88][0]	= 8'h03;
		inst_bytes	[88][1]	= 8'h81;
		inst_bytes	[88][2]	= 8'h01;
		inst_bytes	[88][3]	= 8'h02;
		inst_bytes	[88][4]	= 8'h03;
		inst_bytes	[88][5]	= 8'h04;
		inst_size	[88]		= 4'd6;

		inst_bytes	[89][0]	= 8'h03;
		inst_bytes	[89][1]	= 8'h84;
		inst_bytes	[89][2]	= 8'h52;
		inst_bytes	[89][3]	= 8'h01;
		inst_bytes	[89][4]	= 8'h02;
		inst_bytes	[89][5]	= 8'h03;
		inst_bytes	[89][6]	= 8'h04;
		inst_size	[89]		= 4'd7;

		inst_bytes	[90][0]	= 8'h03;
		inst_bytes	[90][1]	= 8'hC1;
		inst_size	[90]		= 4'd2;

		inst_bytes	[91][0]	= 8'h24;
		inst_bytes	[91][1]	= 8'h11;
		inst_size	[91]		= 4'd2;

		inst_bytes	[92][0]	= 8'h66;
		inst_bytes	[92][1]	= 8'h25;
		inst_bytes	[92][2]	= 8'h11;
		inst_bytes	[92][3]	= 8'h12;
		inst_size	[92]		= 4'd4;

		inst_bytes	[93][0]	= 8'h25;
		inst_bytes	[93][1]	= 8'h11;
		inst_bytes	[93][2]	= 8'h12;
		inst_bytes	[93][3]	= 8'h13;
		inst_bytes	[93][4]	= 8'h14;
		inst_size	[93]		= 4'd5;

		inst_bytes	[94][0]	= 8'h80;
		inst_bytes	[94][1]	= 8'h21;
		inst_bytes	[94][2]	= 8'h11;
		inst_size	[94]		= 4'd3;

		inst_bytes	[95][0]	= 8'h80;
		inst_bytes	[95][1]	= 8'h24;
		inst_bytes	[95][2]	= 8'h52;
		inst_bytes	[95][3]	= 8'h11;
		inst_size	[95]		= 4'd4;

		inst_bytes	[96][0]	= 8'h80;
		inst_bytes	[96][1]	= 8'h25;
		inst_bytes	[96][2]	= 8'h01;
		inst_bytes	[96][3]	= 8'h02;
		inst_bytes	[96][4]	= 8'h03;
		inst_bytes	[96][5]	= 8'h04;
		inst_bytes	[96][6]	= 8'h11;
		inst_size	[96]		= 4'd7;

		inst_bytes	[97][0]	= 8'h80;
		inst_bytes	[97][1]	= 8'h61;
		inst_bytes	[97][2]	= 8'h01;
		inst_bytes	[97][3]	= 8'h11;
		inst_size	[97]		= 4'd4;

		inst_bytes	[98][0]	= 8'h80;
		inst_bytes	[98][1]	= 8'h64;
		inst_bytes	[98][2]	= 8'h52;
		inst_bytes	[98][3]	= 8'h01;
		inst_bytes	[98][4]	= 8'h11;
		inst_size	[98]		= 4'd5;

		inst_bytes	[99][0]	= 8'h80;
		inst_bytes	[99][1]	= 8'hA1;
		inst_bytes	[99][2]	= 8'h01;
		inst_bytes	[99][3]	= 8'h02;
		inst_bytes	[99][4]	= 8'h03;
		inst_bytes	[99][5]	= 8'h04;
		inst_bytes	[99][6]	= 8'h11;
		inst_size	[99]		= 4'd7;

		inst_bytes	[100][0]	= 8'h80;
		inst_bytes	[100][1]	= 8'hA4;
		inst_bytes	[100][2]	= 8'h52;
		inst_bytes	[100][3]	= 8'h01;
		inst_bytes	[100][4]	= 8'h02;
		inst_bytes	[100][5]	= 8'h03;
		inst_bytes	[100][6]	= 8'h04;
		inst_bytes	[100][7]	= 8'h11;
		inst_size	[100]		= 4'd8;

		inst_bytes	[101][0]	= 8'h80;
		inst_bytes	[101][1]	= 8'hE1;
		inst_bytes	[101][2]	= 8'h11;
		inst_size	[101]		= 4'd3;

		inst_bytes	[102][0]	= 8'h66;
		inst_bytes	[102][1]	= 8'h81;
		inst_bytes	[102][2]	= 8'h21;
		inst_bytes	[102][3]	= 8'h11;
		inst_bytes	[102][4]	= 8'h12;
		inst_size	[102]		= 4'd5;

		inst_bytes	[103][0]	= 8'h66;
		inst_bytes	[103][1]	= 8'h81;
		inst_bytes	[103][2]	= 8'h24;
		inst_bytes	[103][3]	= 8'h52;
		inst_bytes	[103][4]	= 8'h11;
		inst_bytes	[103][5]	= 8'h12;
		inst_size	[103]		= 4'd6;

		inst_bytes	[104][0]	= 8'h66;
		inst_bytes	[104][1]	= 8'h81;
		inst_bytes	[104][2]	= 8'h25;
		inst_bytes	[104][3]	= 8'h01;
		inst_bytes	[104][4]	= 8'h02;
		inst_bytes	[104][5]	= 8'h03;
		inst_bytes	[104][6]	= 8'h04;
		inst_bytes	[104][7]	= 8'h11;
		inst_bytes	[104][8]	= 8'h12;
		inst_size	[104]		= 4'd9;

		inst_bytes	[105][0]	= 8'h66;
		inst_bytes	[105][1]	= 8'h81;
		inst_bytes	[105][2]	= 8'h61;
		inst_bytes	[105][3]	= 8'h01;
		inst_bytes	[105][4]	= 8'h11;
		inst_bytes	[105][5]	= 8'h12;
		inst_size	[105]		= 4'd6;

		inst_bytes	[106][0]	= 8'h66;
		inst_bytes	[106][1]	= 8'h81;
		inst_bytes	[106][2]	= 8'h64;
		inst_bytes	[106][3]	= 8'h52;
		inst_bytes	[106][4]	= 8'h01;
		inst_bytes	[106][5]	= 8'h11;
		inst_bytes	[106][6]	= 8'h12;
		inst_size	[106]		= 4'd7;

		inst_bytes	[107][0]	= 8'h66;
		inst_bytes	[107][1]	= 8'h81;
		inst_bytes	[107][2]	= 8'hA1;
		inst_bytes	[107][3]	= 8'h01;
		inst_bytes	[107][4]	= 8'h02;
		inst_bytes	[107][5]	= 8'h03;
		inst_bytes	[107][6]	= 8'h04;
		inst_bytes	[107][7]	= 8'h11;
		inst_bytes	[107][8]	= 8'h12;
		inst_size	[107]		= 4'd9;

		inst_bytes	[108][0]	= 8'h66;
		inst_bytes	[108][1]	= 8'h81;
		inst_bytes	[108][2]	= 8'hA4;
		inst_bytes	[108][3]	= 8'h52;
		inst_bytes	[108][4]	= 8'h01;
		inst_bytes	[108][5]	= 8'h02;
		inst_bytes	[108][6]	= 8'h03;
		inst_bytes	[108][7]	= 8'h04;
		inst_bytes	[108][8]	= 8'h11;
		inst_bytes	[108][9]	= 8'h12;
		inst_size	[108]		= 4'd10;

		inst_bytes	[109][0]	= 8'h66;
		inst_bytes	[109][1]	= 8'h81;
		inst_bytes	[109][2]	= 8'hE1;
		inst_bytes	[109][3]	= 8'h11;
		inst_bytes	[109][4]	= 8'h12;
		inst_size	[109]		= 4'd5;

		inst_bytes	[110][0]	= 8'h81;
		inst_bytes	[110][1]	= 8'h21;
		inst_bytes	[110][2]	= 8'h11;
		inst_bytes	[110][3]	= 8'h12;
		inst_bytes	[110][4]	= 8'h13;
		inst_bytes	[110][5]	= 8'h14;
		inst_size	[110]		= 4'd6;

		inst_bytes	[111][0]	= 8'h81;
		inst_bytes	[111][1]	= 8'h24;
		inst_bytes	[111][2]	= 8'h52;
		inst_bytes	[111][3]	= 8'h11;
		inst_bytes	[111][4]	= 8'h12;
		inst_bytes	[111][5]	= 8'h13;
		inst_bytes	[111][6]	= 8'h14;
		inst_size	[111]		= 4'd7;

		inst_bytes	[112][0]	= 8'h81;
		inst_bytes	[112][1]	= 8'h25;
		inst_bytes	[112][2]	= 8'h01;
		inst_bytes	[112][3]	= 8'h02;
		inst_bytes	[112][4]	= 8'h03;
		inst_bytes	[112][5]	= 8'h04;
		inst_bytes	[112][6]	= 8'h11;
		inst_bytes	[112][7]	= 8'h12;
		inst_bytes	[112][8]	= 8'h13;
		inst_bytes	[112][9]	= 8'h14;
		inst_size	[112]		= 4'd10;

		inst_bytes	[113][0]	= 8'h81;
		inst_bytes	[113][1]	= 8'h61;
		inst_bytes	[113][2]	= 8'h01;
		inst_bytes	[113][3]	= 8'h11;
		inst_bytes	[113][4]	= 8'h12;
		inst_bytes	[113][5]	= 8'h13;
		inst_bytes	[113][6]	= 8'h14;
		inst_size	[113]		= 4'd7;

		inst_bytes	[114][0]	= 8'h81;
		inst_bytes	[114][1]	= 8'h64;
		inst_bytes	[114][2]	= 8'h52;
		inst_bytes	[114][3]	= 8'h01;
		inst_bytes	[114][4]	= 8'h11;
		inst_bytes	[114][5]	= 8'h12;
		inst_bytes	[114][6]	= 8'h13;
		inst_bytes	[114][7]	= 8'h14;
		inst_size	[114]		= 4'd8;

		inst_bytes	[115][0]	= 8'h81;
		inst_bytes	[115][1]	= 8'hA1;
		inst_bytes	[115][2]	= 8'h01;
		inst_bytes	[115][3]	= 8'h02;
		inst_bytes	[115][4]	= 8'h03;
		inst_bytes	[115][5]	= 8'h04;
		inst_bytes	[115][6]	= 8'h11;
		inst_bytes	[115][7]	= 8'h12;
		inst_bytes	[115][8]	= 8'h13;
		inst_bytes	[115][9]	= 8'h14;
		inst_size	[115]		= 4'd10;

		inst_bytes	[116][0]	= 8'h81;
		inst_bytes	[116][1]	= 8'hA4;
		inst_bytes	[116][2]	= 8'h52;
		inst_bytes	[116][3]	= 8'h01;
		inst_bytes	[116][4]	= 8'h02;
		inst_bytes	[116][5]	= 8'h03;
		inst_bytes	[116][6]	= 8'h04;
		inst_bytes	[116][7]	= 8'h11;
		inst_bytes	[116][8]	= 8'h12;
		inst_bytes	[116][9]	= 8'h13;
		inst_bytes	[116][10]	= 8'h14;
		inst_size	[116]		= 4'd11;

		inst_bytes	[117][0]	= 8'h81;
		inst_bytes	[117][1]	= 8'hE1;
		inst_bytes	[117][2]	= 8'h11;
		inst_bytes	[117][3]	= 8'h12;
		inst_bytes	[117][4]	= 8'h13;
		inst_bytes	[117][5]	= 8'h14;
		inst_size	[117]		= 4'd6;

		inst_bytes	[118][0]	= 8'h83;
		inst_bytes	[118][1]	= 8'h21;
		inst_bytes	[118][2]	= 8'h11;
		inst_size	[118]		= 4'd3;

		inst_bytes	[119][0]	= 8'h83;
		inst_bytes	[119][1]	= 8'h24;
		inst_bytes	[119][2]	= 8'h52;
		inst_bytes	[119][3]	= 8'h11;
		inst_size	[119]		= 4'd4;

		inst_bytes	[120][0]	= 8'h83;
		inst_bytes	[120][1]	= 8'h25;
		inst_bytes	[120][2]	= 8'h01;
		inst_bytes	[120][3]	= 8'h02;
		inst_bytes	[120][4]	= 8'h03;
		inst_bytes	[120][5]	= 8'h04;
		inst_bytes	[120][6]	= 8'h11;
		inst_size	[120]		= 4'd7;

		inst_bytes	[121][0]	= 8'h83;
		inst_bytes	[121][1]	= 8'h61;
		inst_bytes	[121][2]	= 8'h01;
		inst_bytes	[121][3]	= 8'h11;
		inst_size	[121]		= 4'd4;

		inst_bytes	[122][0]	= 8'h83;
		inst_bytes	[122][1]	= 8'h64;
		inst_bytes	[122][2]	= 8'h52;
		inst_bytes	[122][3]	= 8'h01;
		inst_bytes	[122][4]	= 8'h11;
		inst_size	[122]		= 4'd5;

		inst_bytes	[123][0]	= 8'h83;
		inst_bytes	[123][1]	= 8'hA1;
		inst_bytes	[123][2]	= 8'h01;
		inst_bytes	[123][3]	= 8'h02;
		inst_bytes	[123][4]	= 8'h03;
		inst_bytes	[123][5]	= 8'h04;
		inst_bytes	[123][6]	= 8'h11;
		inst_size	[123]		= 4'd7;

		inst_bytes	[124][0]	= 8'h83;
		inst_bytes	[124][1]	= 8'hA4;
		inst_bytes	[124][2]	= 8'h52;
		inst_bytes	[124][3]	= 8'h01;
		inst_bytes	[124][4]	= 8'h02;
		inst_bytes	[124][5]	= 8'h03;
		inst_bytes	[124][6]	= 8'h04;
		inst_bytes	[124][7]	= 8'h11;
		inst_size	[124]		= 4'd8;

		inst_bytes	[125][0]	= 8'h83;
		inst_bytes	[125][1]	= 8'hE1;
		inst_bytes	[125][2]	= 8'h11;
		inst_size	[125]		= 4'd3;

		inst_bytes	[126][0]	= 8'h83;
		inst_bytes	[126][1]	= 8'h21;
		inst_bytes	[126][2]	= 8'h11;
		inst_size	[126]		= 4'd3;

		inst_bytes	[127][0]	= 8'h83;
		inst_bytes	[127][1]	= 8'h24;
		inst_bytes	[127][2]	= 8'h52;
		inst_bytes	[127][3]	= 8'h11;
		inst_size	[127]		= 4'd4;

		inst_bytes	[128][0]	= 8'h83;
		inst_bytes	[128][1]	= 8'h25;
		inst_bytes	[128][2]	= 8'h01;
		inst_bytes	[128][3]	= 8'h02;
		inst_bytes	[128][4]	= 8'h03;
		inst_bytes	[128][5]	= 8'h04;
		inst_bytes	[128][6]	= 8'h11;
		inst_size	[128]		= 4'd7;

		inst_bytes	[129][0]	= 8'h83;
		inst_bytes	[129][1]	= 8'h61;
		inst_bytes	[129][2]	= 8'h01;
		inst_bytes	[129][3]	= 8'h11;
		inst_size	[129]		= 4'd4;

		inst_bytes	[130][0]	= 8'h83;
		inst_bytes	[130][1]	= 8'h64;
		inst_bytes	[130][2]	= 8'h52;
		inst_bytes	[130][3]	= 8'h01;
		inst_bytes	[130][4]	= 8'h11;
		inst_size	[130]		= 4'd5;

		inst_bytes	[131][0]	= 8'h83;
		inst_bytes	[131][1]	= 8'hA1;
		inst_bytes	[131][2]	= 8'h01;
		inst_bytes	[131][3]	= 8'h02;
		inst_bytes	[131][4]	= 8'h03;
		inst_bytes	[131][5]	= 8'h04;
		inst_bytes	[131][6]	= 8'h11;
		inst_size	[131]		= 4'd7;

		inst_bytes	[132][0]	= 8'h83;
		inst_bytes	[132][1]	= 8'hA4;
		inst_bytes	[132][2]	= 8'h52;
		inst_bytes	[132][3]	= 8'h01;
		inst_bytes	[132][4]	= 8'h02;
		inst_bytes	[132][5]	= 8'h03;
		inst_bytes	[132][6]	= 8'h04;
		inst_bytes	[132][7]	= 8'h11;
		inst_size	[132]		= 4'd8;

		inst_bytes	[133][0]	= 8'h83;
		inst_bytes	[133][1]	= 8'hE1;
		inst_bytes	[133][2]	= 8'h11;
		inst_size	[133]		= 4'd3;

		inst_bytes	[134][0]	= 8'h20;
		inst_bytes	[134][1]	= 8'h01;
		inst_size	[134]		= 4'd2;

		inst_bytes	[135][0]	= 8'h20;
		inst_bytes	[135][1]	= 8'h04;
		inst_bytes	[135][2]	= 8'h52;
		inst_size	[135]		= 4'd3;

		inst_bytes	[136][0]	= 8'h20;
		inst_bytes	[136][1]	= 8'h05;
		inst_bytes	[136][2]	= 8'h01;
		inst_bytes	[136][3]	= 8'h02;
		inst_bytes	[136][4]	= 8'h03;
		inst_bytes	[136][5]	= 8'h04;
		inst_size	[136]		= 4'd6;

		inst_bytes	[137][0]	= 8'h20;
		inst_bytes	[137][1]	= 8'h41;
		inst_bytes	[137][2]	= 8'h01;
		inst_size	[137]		= 4'd3;

		inst_bytes	[138][0]	= 8'h20;
		inst_bytes	[138][1]	= 8'h44;
		inst_bytes	[138][2]	= 8'h52;
		inst_bytes	[138][3]	= 8'h01;
		inst_size	[138]		= 4'd4;

		inst_bytes	[139][0]	= 8'h20;
		inst_bytes	[139][1]	= 8'h81;
		inst_bytes	[139][2]	= 8'h01;
		inst_bytes	[139][3]	= 8'h02;
		inst_bytes	[139][4]	= 8'h03;
		inst_bytes	[139][5]	= 8'h04;
		inst_size	[139]		= 4'd6;

		inst_bytes	[140][0]	= 8'h20;
		inst_bytes	[140][1]	= 8'h84;
		inst_bytes	[140][2]	= 8'h52;
		inst_bytes	[140][3]	= 8'h01;
		inst_bytes	[140][4]	= 8'h02;
		inst_bytes	[140][5]	= 8'h03;
		inst_bytes	[140][6]	= 8'h04;
		inst_size	[140]		= 4'd7;

		inst_bytes	[141][0]	= 8'h20;
		inst_bytes	[141][1]	= 8'hC1;
		inst_size	[141]		= 4'd2;

		inst_bytes	[142][0]	= 8'h21;
		inst_bytes	[142][1]	= 8'h01;
		inst_size	[142]		= 4'd2;

		inst_bytes	[143][0]	= 8'h21;
		inst_bytes	[143][1]	= 8'h04;
		inst_bytes	[143][2]	= 8'h52;
		inst_size	[143]		= 4'd3;

		inst_bytes	[144][0]	= 8'h21;
		inst_bytes	[144][1]	= 8'h05;
		inst_bytes	[144][2]	= 8'h01;
		inst_bytes	[144][3]	= 8'h02;
		inst_bytes	[144][4]	= 8'h03;
		inst_bytes	[144][5]	= 8'h04;
		inst_size	[144]		= 4'd6;

		inst_bytes	[145][0]	= 8'h21;
		inst_bytes	[145][1]	= 8'h41;
		inst_bytes	[145][2]	= 8'h01;
		inst_size	[145]		= 4'd3;

		inst_bytes	[146][0]	= 8'h21;
		inst_bytes	[146][1]	= 8'h44;
		inst_bytes	[146][2]	= 8'h52;
		inst_bytes	[146][3]	= 8'h01;
		inst_size	[146]		= 4'd4;

		inst_bytes	[147][0]	= 8'h21;
		inst_bytes	[147][1]	= 8'h81;
		inst_bytes	[147][2]	= 8'h01;
		inst_bytes	[147][3]	= 8'h02;
		inst_bytes	[147][4]	= 8'h03;
		inst_bytes	[147][5]	= 8'h04;
		inst_size	[147]		= 4'd6;

		inst_bytes	[148][0]	= 8'h21;
		inst_bytes	[148][1]	= 8'h84;
		inst_bytes	[148][2]	= 8'h52;
		inst_bytes	[148][3]	= 8'h01;
		inst_bytes	[148][4]	= 8'h02;
		inst_bytes	[148][5]	= 8'h03;
		inst_bytes	[148][6]	= 8'h04;
		inst_size	[148]		= 4'd7;

		inst_bytes	[149][0]	= 8'h21;
		inst_bytes	[149][1]	= 8'hC1;
		inst_size	[149]		= 4'd2;

		inst_bytes	[150][0]	= 8'h21;
		inst_bytes	[150][1]	= 8'h01;
		inst_size	[150]		= 4'd2;

		inst_bytes	[151][0]	= 8'h21;
		inst_bytes	[151][1]	= 8'h04;
		inst_bytes	[151][2]	= 8'h52;
		inst_size	[151]		= 4'd3;

		inst_bytes	[152][0]	= 8'h21;
		inst_bytes	[152][1]	= 8'h05;
		inst_bytes	[152][2]	= 8'h01;
		inst_bytes	[152][3]	= 8'h02;
		inst_bytes	[152][4]	= 8'h03;
		inst_bytes	[152][5]	= 8'h04;
		inst_size	[152]		= 4'd6;

		inst_bytes	[153][0]	= 8'h21;
		inst_bytes	[153][1]	= 8'h41;
		inst_bytes	[153][2]	= 8'h01;
		inst_size	[153]		= 4'd3;

		inst_bytes	[154][0]	= 8'h21;
		inst_bytes	[154][1]	= 8'h44;
		inst_bytes	[154][2]	= 8'h52;
		inst_bytes	[154][3]	= 8'h01;
		inst_size	[154]		= 4'd4;

		inst_bytes	[155][0]	= 8'h21;
		inst_bytes	[155][1]	= 8'h81;
		inst_bytes	[155][2]	= 8'h01;
		inst_bytes	[155][3]	= 8'h02;
		inst_bytes	[155][4]	= 8'h03;
		inst_bytes	[155][5]	= 8'h04;
		inst_size	[155]		= 4'd6;

		inst_bytes	[156][0]	= 8'h21;
		inst_bytes	[156][1]	= 8'h84;
		inst_bytes	[156][2]	= 8'h52;
		inst_bytes	[156][3]	= 8'h01;
		inst_bytes	[156][4]	= 8'h02;
		inst_bytes	[156][5]	= 8'h03;
		inst_bytes	[156][6]	= 8'h04;
		inst_size	[156]		= 4'd7;

		inst_bytes	[157][0]	= 8'h21;
		inst_bytes	[157][1]	= 8'hC1;
		inst_size	[157]		= 4'd2;

		inst_bytes	[158][0]	= 8'h22;
		inst_bytes	[158][1]	= 8'h01;
		inst_size	[158]		= 4'd2;

		inst_bytes	[159][0]	= 8'h22;
		inst_bytes	[159][1]	= 8'h04;
		inst_bytes	[159][2]	= 8'h52;
		inst_size	[159]		= 4'd3;

		inst_bytes	[160][0]	= 8'h22;
		inst_bytes	[160][1]	= 8'h05;
		inst_bytes	[160][2]	= 8'h01;
		inst_bytes	[160][3]	= 8'h02;
		inst_bytes	[160][4]	= 8'h03;
		inst_bytes	[160][5]	= 8'h04;
		inst_size	[160]		= 4'd6;

		inst_bytes	[161][0]	= 8'h22;
		inst_bytes	[161][1]	= 8'h41;
		inst_bytes	[161][2]	= 8'h01;
		inst_size	[161]		= 4'd3;

		inst_bytes	[162][0]	= 8'h22;
		inst_bytes	[162][1]	= 8'h44;
		inst_bytes	[162][2]	= 8'h52;
		inst_bytes	[162][3]	= 8'h01;
		inst_size	[162]		= 4'd4;

		inst_bytes	[163][0]	= 8'h22;
		inst_bytes	[163][1]	= 8'h81;
		inst_bytes	[163][2]	= 8'h01;
		inst_bytes	[163][3]	= 8'h02;
		inst_bytes	[163][4]	= 8'h03;
		inst_bytes	[163][5]	= 8'h04;
		inst_size	[163]		= 4'd6;

		inst_bytes	[164][0]	= 8'h22;
		inst_bytes	[164][1]	= 8'h84;
		inst_bytes	[164][2]	= 8'h52;
		inst_bytes	[164][3]	= 8'h01;
		inst_bytes	[164][4]	= 8'h02;
		inst_bytes	[164][5]	= 8'h03;
		inst_bytes	[164][6]	= 8'h04;
		inst_size	[164]		= 4'd7;

		inst_bytes	[165][0]	= 8'h22;
		inst_bytes	[165][1]	= 8'hC1;
		inst_size	[165]		= 4'd2;

		inst_bytes	[166][0]	= 8'h23;
		inst_bytes	[166][1]	= 8'h01;
		inst_size	[166]		= 4'd2;

		inst_bytes	[167][0]	= 8'h23;
		inst_bytes	[167][1]	= 8'h04;
		inst_bytes	[167][2]	= 8'h52;
		inst_size	[167]		= 4'd3;

		inst_bytes	[168][0]	= 8'h23;
		inst_bytes	[168][1]	= 8'h05;
		inst_bytes	[168][2]	= 8'h01;
		inst_bytes	[168][3]	= 8'h02;
		inst_bytes	[168][4]	= 8'h03;
		inst_bytes	[168][5]	= 8'h04;
		inst_size	[168]		= 4'd6;

		inst_bytes	[169][0]	= 8'h23;
		inst_bytes	[169][1]	= 8'h41;
		inst_bytes	[169][2]	= 8'h01;
		inst_size	[169]		= 4'd3;

		inst_bytes	[170][0]	= 8'h23;
		inst_bytes	[170][1]	= 8'h44;
		inst_bytes	[170][2]	= 8'h52;
		inst_bytes	[170][3]	= 8'h01;
		inst_size	[170]		= 4'd4;

		inst_bytes	[171][0]	= 8'h23;
		inst_bytes	[171][1]	= 8'h81;
		inst_bytes	[171][2]	= 8'h01;
		inst_bytes	[171][3]	= 8'h02;
		inst_bytes	[171][4]	= 8'h03;
		inst_bytes	[171][5]	= 8'h04;
		inst_size	[171]		= 4'd6;

		inst_bytes	[172][0]	= 8'h23;
		inst_bytes	[172][1]	= 8'h84;
		inst_bytes	[172][2]	= 8'h52;
		inst_bytes	[172][3]	= 8'h01;
		inst_bytes	[172][4]	= 8'h02;
		inst_bytes	[172][5]	= 8'h03;
		inst_bytes	[172][6]	= 8'h04;
		inst_size	[172]		= 4'd7;

		inst_bytes	[173][0]	= 8'h23;
		inst_bytes	[173][1]	= 8'hC1;
		inst_size	[173]		= 4'd2;

		inst_bytes	[174][0]	= 8'h23;
		inst_bytes	[174][1]	= 8'h01;
		inst_size	[174]		= 4'd2;

		inst_bytes	[175][0]	= 8'h23;
		inst_bytes	[175][1]	= 8'h04;
		inst_bytes	[175][2]	= 8'h52;
		inst_size	[175]		= 4'd3;

		inst_bytes	[176][0]	= 8'h23;
		inst_bytes	[176][1]	= 8'h05;
		inst_bytes	[176][2]	= 8'h01;
		inst_bytes	[176][3]	= 8'h02;
		inst_bytes	[176][4]	= 8'h03;
		inst_bytes	[176][5]	= 8'h04;
		inst_size	[176]		= 4'd6;

		inst_bytes	[177][0]	= 8'h23;
		inst_bytes	[177][1]	= 8'h41;
		inst_bytes	[177][2]	= 8'h01;
		inst_size	[177]		= 4'd3;

		inst_bytes	[178][0]	= 8'h23;
		inst_bytes	[178][1]	= 8'h44;
		inst_bytes	[178][2]	= 8'h52;
		inst_bytes	[178][3]	= 8'h01;
		inst_size	[178]		= 4'd4;

		inst_bytes	[179][0]	= 8'h23;
		inst_bytes	[179][1]	= 8'h81;
		inst_bytes	[179][2]	= 8'h01;
		inst_bytes	[179][3]	= 8'h02;
		inst_bytes	[179][4]	= 8'h03;
		inst_bytes	[179][5]	= 8'h04;
		inst_size	[179]		= 4'd6;

		inst_bytes	[180][0]	= 8'h23;
		inst_bytes	[180][1]	= 8'h84;
		inst_bytes	[180][2]	= 8'h52;
		inst_bytes	[180][3]	= 8'h01;
		inst_bytes	[180][4]	= 8'h02;
		inst_bytes	[180][5]	= 8'h03;
		inst_bytes	[180][6]	= 8'h04;
		inst_size	[180]		= 4'd7;

		inst_bytes	[181][0]	= 8'h23;
		inst_bytes	[181][1]	= 8'hC1;
		inst_size	[181]		= 4'd2;

		inst_bytes	[182][0]	= 8'h66;
		inst_bytes	[182][1]	= 8'hE8;
		inst_bytes	[182][2]	= 8'h11;
		inst_bytes	[182][3]	= 8'h12;
		inst_size	[182]		= 4'd4;

		inst_bytes	[183][0]	= 8'hE8;
		inst_bytes	[183][1]	= 8'h11;
		inst_bytes	[183][2]	= 8'h12;
		inst_bytes	[183][3]	= 8'h13;
		inst_bytes	[183][4]	= 8'h14;
		inst_size	[183]		= 4'd5;

		inst_bytes	[184][0]	= 8'hFF;
		inst_bytes	[184][1]	= 8'h11;
		inst_size	[184]		= 4'd2;

		inst_bytes	[185][0]	= 8'hFF;
		inst_bytes	[185][1]	= 8'h14;
		inst_bytes	[185][2]	= 8'h52;
		inst_size	[185]		= 4'd3;

		inst_bytes	[186][0]	= 8'hFF;
		inst_bytes	[186][1]	= 8'h15;
		inst_bytes	[186][2]	= 8'h01;
		inst_bytes	[186][3]	= 8'h02;
		inst_bytes	[186][4]	= 8'h03;
		inst_bytes	[186][5]	= 8'h04;
		inst_size	[186]		= 4'd6;

		inst_bytes	[187][0]	= 8'hFF;
		inst_bytes	[187][1]	= 8'h51;
		inst_bytes	[187][2]	= 8'h01;
		inst_size	[187]		= 4'd3;

		inst_bytes	[188][0]	= 8'hFF;
		inst_bytes	[188][1]	= 8'h54;
		inst_bytes	[188][2]	= 8'h52;
		inst_bytes	[188][3]	= 8'h01;
		inst_size	[188]		= 4'd4;

		inst_bytes	[189][0]	= 8'hFF;
		inst_bytes	[189][1]	= 8'h91;
		inst_bytes	[189][2]	= 8'h01;
		inst_bytes	[189][3]	= 8'h02;
		inst_bytes	[189][4]	= 8'h04;
		inst_bytes	[189][5]	= 8'h04;
		inst_size	[189]		= 4'd6;

		inst_bytes	[190][0]	= 8'hFF;
		inst_bytes	[190][1]	= 8'h94;
		inst_bytes	[190][2]	= 8'h52;
		inst_bytes	[190][3]	= 8'h01;
		inst_bytes	[190][4]	= 8'h02;
		inst_bytes	[190][5]	= 8'h03;
		inst_bytes	[190][6]	= 8'h04;
		inst_size	[190]		= 4'd7;

		inst_bytes	[191][0]	= 8'hFF;
		inst_bytes	[191][1]	= 8'hD1;
		inst_size	[191]		= 4'd2;

		inst_bytes	[192][0]	= 8'hFF;
		inst_bytes	[192][1]	= 8'h11;
		inst_size	[192]		= 4'd2;

		inst_bytes	[193][0]	= 8'hFF;
		inst_bytes	[193][1]	= 8'h14;
		inst_bytes	[193][2]	= 8'h52;
		inst_size	[193]		= 4'd3;

		inst_bytes	[194][0]	= 8'hFF;
		inst_bytes	[194][1]	= 8'h15;
		inst_bytes	[194][2]	= 8'h01;
		inst_bytes	[194][3]	= 8'h02;
		inst_bytes	[194][4]	= 8'h03;
		inst_bytes	[194][5]	= 8'h04;
		inst_size	[194]		= 4'd6;

		inst_bytes	[195][0]	= 8'hFF;
		inst_bytes	[195][1]	= 8'h51;
		inst_bytes	[195][2]	= 8'h01;
		inst_size	[195]		= 4'd3;

		inst_bytes	[196][0]	= 8'hFF;
		inst_bytes	[196][1]	= 8'h54;
		inst_bytes	[196][2]	= 8'h52;
		inst_bytes	[196][3]	= 8'h01;
		inst_size	[196]		= 4'd4;

		inst_bytes	[197][0]	= 8'hFF;
		inst_bytes	[197][1]	= 8'h91;
		inst_bytes	[197][2]	= 8'h01;
		inst_bytes	[197][3]	= 8'h02;
		inst_bytes	[197][4]	= 8'h04;
		inst_bytes	[197][5]	= 8'h04;
		inst_size	[197]		= 4'd6;

		inst_bytes	[198][0]	= 8'hFF;
		inst_bytes	[198][1]	= 8'h94;
		inst_bytes	[198][2]	= 8'h52;
		inst_bytes	[198][3]	= 8'h01;
		inst_bytes	[198][4]	= 8'h02;
		inst_bytes	[198][5]	= 8'h03;
		inst_bytes	[198][6]	= 8'h04;
		inst_size	[198]		= 4'd7;

		inst_bytes	[199][0]	= 8'hFF;
		inst_bytes	[199][1]	= 8'hD1;
		inst_size	[199]		= 4'd2;

		inst_bytes	[200][0]	= 8'h9A;
		inst_bytes	[200][1]	= 8'h0F;
		inst_bytes	[200][2]	= 8'h10;
		inst_bytes	[200][3]	= 8'h11;
		inst_bytes	[200][4]	= 8'h12;
		inst_bytes	[200][5]	= 8'h13;
		inst_bytes	[200][6]	= 8'h14;
		inst_size	[200]		= 4'd7;

		inst_bytes	[201][0]	= 8'hFC;
		inst_size	[201]		= 4'd1;

		inst_bytes	[202][0]	= 8'h0F;
		inst_bytes	[202][1]	= 8'h42;
		inst_bytes	[202][2]	= 8'h01;
		inst_size	[202]		= 4'd3;

		inst_bytes	[203][0]	= 8'h0F;
		inst_bytes	[203][1]	= 8'h42;
		inst_bytes	[203][2]	= 8'h04;
		inst_bytes	[203][3]	= 8'h52;
		inst_size	[203]		= 4'd4;

		inst_bytes	[204][0]	= 8'h0F;
		inst_bytes	[204][1]	= 8'h42;
		inst_bytes	[204][2]	= 8'h05;
		inst_bytes	[204][3]	= 8'h01;
		inst_bytes	[204][4]	= 8'h02;
		inst_bytes	[204][5]	= 8'h03;
		inst_bytes	[204][6]	= 8'h04;
		inst_size	[204]		= 4'd7;

		inst_bytes	[205][0]	= 8'h0F;
		inst_bytes	[205][1]	= 8'h42;
		inst_bytes	[205][2]	= 8'h41;
		inst_bytes	[205][3]	= 8'h01;
		inst_size	[205]		= 4'd4;

		inst_bytes	[206][0]	= 8'h0F;
		inst_bytes	[206][1]	= 8'h42;
		inst_bytes	[206][2]	= 8'h44;
		inst_bytes	[206][3]	= 8'h52;
		inst_bytes	[206][4]	= 8'h01;
		inst_size	[206]		= 4'd5;

		inst_bytes	[207][0]	= 8'h0F;
		inst_bytes	[207][1]	= 8'h42;
		inst_bytes	[207][2]	= 8'h81;
		inst_bytes	[207][3]	= 8'h01;
		inst_bytes	[207][4]	= 8'h02;
		inst_bytes	[207][5]	= 8'h03;
		inst_bytes	[207][6]	= 8'h04;
		inst_size	[207]		= 4'd7;

		inst_bytes	[208][0]	= 8'h0F;
		inst_bytes	[208][1]	= 8'h42;
		inst_bytes	[208][2]	= 8'h84;
		inst_bytes	[208][3]	= 8'h52;
		inst_bytes	[208][4]	= 8'h01;
		inst_bytes	[208][5]	= 8'h02;
		inst_bytes	[208][6]	= 8'h03;
		inst_bytes	[208][7]	= 8'h04;
		inst_size	[208]		= 4'd8;

		inst_bytes	[209][0]	= 8'h0F;
		inst_bytes	[209][1]	= 8'h42;
		inst_bytes	[209][2]	= 8'hC1;
		inst_size	[209]		= 4'd3;

		inst_bytes	[210][0]	= 8'h0F;
		inst_bytes	[210][1]	= 8'h42;
		inst_bytes	[210][2]	= 8'h01;
		inst_size	[210]		= 4'd3;

		inst_bytes	[211][0]	= 8'h0F;
		inst_bytes	[211][1]	= 8'h42;
		inst_bytes	[211][2]	= 8'h04;
		inst_bytes	[211][3]	= 8'h52;
		inst_size	[211]		= 4'd4;

		inst_bytes	[212][0]	= 8'h0F;
		inst_bytes	[212][1]	= 8'h42;
		inst_bytes	[212][2]	= 8'h05;
		inst_bytes	[212][3]	= 8'h01;
		inst_bytes	[212][4]	= 8'h02;
		inst_bytes	[212][5]	= 8'h03;
		inst_bytes	[212][6]	= 8'h04;
		inst_size	[212]		= 4'd7;

		inst_bytes	[213][0]	= 8'h0F;
		inst_bytes	[213][1]	= 8'h42;
		inst_bytes	[213][2]	= 8'h41;
		inst_bytes	[213][3]	= 8'h01;
		inst_size	[213]		= 4'd4;

		inst_bytes	[214][0]	= 8'h0F;
		inst_bytes	[214][1]	= 8'h42;
		inst_bytes	[214][2]	= 8'h44;
		inst_bytes	[214][3]	= 8'h52;
		inst_bytes	[214][4]	= 8'h01;
		inst_size	[214]		= 4'd5;

		inst_bytes	[215][0]	= 8'h0F;
		inst_bytes	[215][1]	= 8'h42;
		inst_bytes	[215][2]	= 8'h81;
		inst_bytes	[215][3]	= 8'h01;
		inst_bytes	[215][4]	= 8'h02;
		inst_bytes	[215][5]	= 8'h03;
		inst_bytes	[215][6]	= 8'h04;
		inst_size	[215]		= 4'd7;

		inst_bytes	[216][0]	= 8'h0F;
		inst_bytes	[216][1]	= 8'h42;
		inst_bytes	[216][2]	= 8'h84;
		inst_bytes	[216][3]	= 8'h52;
		inst_bytes	[216][4]	= 8'h01;
		inst_bytes	[216][5]	= 8'h02;
		inst_bytes	[216][6]	= 8'h03;
		inst_bytes	[216][7]	= 8'h04;
		inst_size	[216]		= 4'd8;

		inst_bytes	[217][0]	= 8'h0F;
		inst_bytes	[217][1]	= 8'h42;
		inst_bytes	[217][2]	= 8'hC1;
		inst_size	[217]		= 4'd3;

		inst_bytes	[218][0]	= 8'h0F;
		inst_bytes	[218][1]	= 8'hB0;
		inst_bytes	[218][2]	= 8'h01;
		inst_size	[218]		= 4'd3;

		inst_bytes	[219][0]	= 8'h0F;
		inst_bytes	[219][1]	= 8'hB0;
		inst_bytes	[219][2]	= 8'h04;
		inst_bytes	[219][3]	= 8'h52;
		inst_size	[219]		= 4'd4;

		inst_bytes	[220][0]	= 8'h0F;
		inst_bytes	[220][1]	= 8'hB0;
		inst_bytes	[220][2]	= 8'h05;
		inst_bytes	[220][3]	= 8'h01;
		inst_bytes	[220][4]	= 8'h02;
		inst_bytes	[220][5]	= 8'h03;
		inst_bytes	[220][6]	= 8'h04;
		inst_size	[220]		= 4'd7;

		inst_bytes	[221][0]	= 8'h0F;
		inst_bytes	[221][1]	= 8'hB0;
		inst_bytes	[221][2]	= 8'h41;
		inst_bytes	[221][3]	= 8'h01;
		inst_size	[221]		= 4'd4;

		inst_bytes	[222][0]	= 8'h0F;
		inst_bytes	[222][1]	= 8'hB0;
		inst_bytes	[222][2]	= 8'h44;
		inst_bytes	[222][3]	= 8'h52;
		inst_bytes	[222][4]	= 8'h01;
		inst_size	[222]		= 4'd5;

		inst_bytes	[223][0]	= 8'h0F;
		inst_bytes	[223][1]	= 8'hB0;
		inst_bytes	[223][2]	= 8'h81;
		inst_bytes	[223][3]	= 8'h01;
		inst_bytes	[223][4]	= 8'h02;
		inst_bytes	[223][5]	= 8'h03;
		inst_bytes	[223][6]	= 8'h04;
		inst_size	[223]		= 4'd7;

		inst_bytes	[224][0]	= 8'h0F;
		inst_bytes	[224][1]	= 8'hB0;
		inst_bytes	[224][2]	= 8'h84;
		inst_bytes	[224][3]	= 8'h52;
		inst_bytes	[224][4]	= 8'h01;
		inst_bytes	[224][5]	= 8'h02;
		inst_bytes	[224][6]	= 8'h03;
		inst_bytes	[224][7]	= 8'h04;
		inst_size	[224]		= 4'd8;

		inst_bytes	[225][0]	= 8'h0F;
		inst_bytes	[225][1]	= 8'hB0;
		inst_bytes	[225][2]	= 8'hC1;
		inst_size	[225]		= 4'd3;

		inst_bytes	[226][0]	= 8'h0F;
		inst_bytes	[226][1]	= 8'hB1;
		inst_bytes	[226][2]	= 8'h01;
		inst_size	[226]		= 4'd3;

		inst_bytes	[227][0]	= 8'h0F;
		inst_bytes	[227][1]	= 8'hB1;
		inst_bytes	[227][2]	= 8'h04;
		inst_bytes	[227][3]	= 8'h52;
		inst_size	[227]		= 4'd4;

		inst_bytes	[228][0]	= 8'h0F;
		inst_bytes	[228][1]	= 8'hB1;
		inst_bytes	[228][2]	= 8'h05;
		inst_bytes	[228][3]	= 8'h01;
		inst_bytes	[228][4]	= 8'h02;
		inst_bytes	[228][5]	= 8'h03;
		inst_bytes	[228][6]	= 8'h04;
		inst_size	[228]		= 4'd7;

		inst_bytes	[229][0]	= 8'h0F;
		inst_bytes	[229][1]	= 8'hB1;
		inst_bytes	[229][2]	= 8'h41;
		inst_bytes	[229][3]	= 8'h01;
		inst_size	[229]		= 4'd4;

		inst_bytes	[230][0]	= 8'h0F;
		inst_bytes	[230][1]	= 8'hB1;
		inst_bytes	[230][2]	= 8'h44;
		inst_bytes	[230][3]	= 8'h52;
		inst_bytes	[230][4]	= 8'h01;
		inst_size	[230]		= 4'd5;

		inst_bytes	[231][0]	= 8'h0F;
		inst_bytes	[231][1]	= 8'hB1;
		inst_bytes	[231][2]	= 8'h81;
		inst_bytes	[231][3]	= 8'h01;
		inst_bytes	[231][4]	= 8'h02;
		inst_bytes	[231][5]	= 8'h03;
		inst_bytes	[231][6]	= 8'h04;
		inst_size	[231]		= 4'd7;

		inst_bytes	[232][0]	= 8'h0F;
		inst_bytes	[232][1]	= 8'hB1;
		inst_bytes	[232][2]	= 8'h84;
		inst_bytes	[232][3]	= 8'h52;
		inst_bytes	[232][4]	= 8'h01;
		inst_bytes	[232][5]	= 8'h02;
		inst_bytes	[232][6]	= 8'h03;
		inst_bytes	[232][7]	= 8'h04;
		inst_size	[232]		= 4'd8;

		inst_bytes	[233][0]	= 8'h0F;
		inst_bytes	[233][1]	= 8'hB1;
		inst_bytes	[233][2]	= 8'hC1;
		inst_size	[233]		= 4'd3;

		inst_bytes	[234][0]	= 8'h0F;
		inst_bytes	[234][1]	= 8'hB1;
		inst_bytes	[234][2]	= 8'h01;
		inst_size	[234]		= 4'd3;

		inst_bytes	[235][0]	= 8'h0F;
		inst_bytes	[235][1]	= 8'hB1;
		inst_bytes	[235][2]	= 8'h04;
		inst_bytes	[235][3]	= 8'h52;
		inst_size	[235]		= 4'd4;

		inst_bytes	[236][0]	= 8'h0F;
		inst_bytes	[236][1]	= 8'hB1;
		inst_bytes	[236][2]	= 8'h05;
		inst_bytes	[236][3]	= 8'h01;
		inst_bytes	[236][4]	= 8'h02;
		inst_bytes	[236][5]	= 8'h03;
		inst_bytes	[236][6]	= 8'h04;
		inst_size	[236]		= 4'd7;

		inst_bytes	[237][0]	= 8'h0F;
		inst_bytes	[237][1]	= 8'hB1;
		inst_bytes	[237][2]	= 8'h41;
		inst_bytes	[237][3]	= 8'h01;
		inst_size	[237]		= 4'd4;

		inst_bytes	[238][0]	= 8'h0F;
		inst_bytes	[238][1]	= 8'hB1;
		inst_bytes	[238][2]	= 8'h44;
		inst_bytes	[238][3]	= 8'h52;
		inst_bytes	[238][4]	= 8'h01;
		inst_size	[238]		= 4'd5;

		inst_bytes	[239][0]	= 8'h0F;
		inst_bytes	[239][1]	= 8'hB1;
		inst_bytes	[239][2]	= 8'h81;
		inst_bytes	[239][3]	= 8'h01;
		inst_bytes	[239][4]	= 8'h02;
		inst_bytes	[239][5]	= 8'h03;
		inst_bytes	[239][6]	= 8'h04;
		inst_size	[239]		= 4'd7;

		inst_bytes	[240][0]	= 8'h0F;
		inst_bytes	[240][1]	= 8'hB1;
		inst_bytes	[240][2]	= 8'h84;
		inst_bytes	[240][3]	= 8'h52;
		inst_bytes	[240][4]	= 8'h01;
		inst_bytes	[240][5]	= 8'h02;
		inst_bytes	[240][6]	= 8'h03;
		inst_bytes	[240][7]	= 8'h04;
		inst_size	[240]		= 4'd8;

		inst_bytes	[241][0]	= 8'h0F;
		inst_bytes	[241][1]	= 8'hB1;
		inst_bytes	[241][2]	= 8'hC1;
		inst_size	[241]		= 4'd3;

		inst_bytes	[242][0]	= 8'h27;
		inst_size	[242]		= 4'd1;

		inst_bytes	[243][0]	= 8'hF4;
		inst_size	[243]		= 4'd1;

		inst_bytes	[244][0]	= 8'hFE;
		inst_bytes	[244][1]	= 8'h01;
		inst_size	[244]		= 4'd2;

		inst_bytes	[245][0]	= 8'hFE;
		inst_bytes	[245][1]	= 8'h04;
		inst_bytes	[245][2]	= 8'h52;
		inst_size	[245]		= 4'd3;

		inst_bytes	[246][0]	= 8'hFE;
		inst_bytes	[246][1]	= 8'h05;
		inst_bytes	[246][2]	= 8'h01;
		inst_bytes	[246][3]	= 8'h02;
		inst_bytes	[246][4]	= 8'h03;
		inst_bytes	[246][5]	= 8'h04;
		inst_size	[246]		= 4'd6;

		inst_bytes	[247][0]	= 8'hFE;
		inst_bytes	[247][1]	= 8'h41;
		inst_bytes	[247][2]	= 8'h01;
		inst_size	[247]		= 4'd3;

		inst_bytes	[248][0]	= 8'hFE;
		inst_bytes	[248][1]	= 8'h44;
		inst_bytes	[248][2]	= 8'h52;
		inst_bytes	[248][3]	= 8'h01;
		inst_size	[248]		= 4'd4;

		inst_bytes	[249][0]	= 8'hFE;
		inst_bytes	[249][1]	= 8'h81;
		inst_bytes	[249][2]	= 8'h01;
		inst_bytes	[249][3]	= 8'h02;
		inst_bytes	[249][4]	= 8'h03;
		inst_bytes	[249][5]	= 8'h04;
		inst_size	[249]		= 4'd6;

		inst_bytes	[250][0]	= 8'hFE;
		inst_bytes	[250][1]	= 8'h84;
		inst_bytes	[250][2]	= 8'h52;
		inst_bytes	[250][3]	= 8'h01;
		inst_bytes	[250][4]	= 8'h02;
		inst_bytes	[250][5]	= 8'h03;
		inst_bytes	[250][6]	= 8'h04;
		inst_size	[250]		= 4'd7;

		inst_bytes	[251][0]	= 8'hFE;
		inst_bytes	[251][1]	= 8'hC1;
		inst_size	[251]		= 4'd2;

		inst_bytes	[252][0]	= 8'hFF;
		inst_bytes	[252][1]	= 8'h01;
		inst_size	[252]		= 4'd2;

		inst_bytes	[253][0]	= 8'hFF;
		inst_bytes	[253][1]	= 8'h04;
		inst_bytes	[253][2]	= 8'h52;
		inst_size	[253]		= 4'd3;

		inst_bytes	[254][0]	= 8'hFF;
		inst_bytes	[254][1]	= 8'h05;
		inst_bytes	[254][2]	= 8'h01;
		inst_bytes	[254][3]	= 8'h02;
		inst_bytes	[254][4]	= 8'h03;
		inst_bytes	[254][5]	= 8'h04;
		inst_size	[254]		= 4'd6;

		inst_bytes	[255][0]	= 8'hFF;
		inst_bytes	[255][1]	= 8'h41;
		inst_bytes	[255][2]	= 8'h01;
		inst_size	[255]		= 4'd3;

		inst_bytes	[256][0]	= 8'hFF;
		inst_bytes	[256][1]	= 8'h44;
		inst_bytes	[256][2]	= 8'h52;
		inst_bytes	[256][3]	= 8'h01;
		inst_size	[256]		= 4'd4;

		inst_bytes	[257][0]	= 8'hFF;
		inst_bytes	[257][1]	= 8'h81;
		inst_bytes	[257][2]	= 8'h01;
		inst_bytes	[257][3]	= 8'h02;
		inst_bytes	[257][4]	= 8'h03;
		inst_bytes	[257][5]	= 8'h04;
		inst_size	[257]		= 4'd6;

		inst_bytes	[258][0]	= 8'hFF;
		inst_bytes	[258][1]	= 8'h84;
		inst_bytes	[258][2]	= 8'h52;
		inst_bytes	[258][3]	= 8'h01;
		inst_bytes	[258][4]	= 8'h02;
		inst_bytes	[258][5]	= 8'h03;
		inst_bytes	[258][6]	= 8'h04;
		inst_size	[258]		= 4'd7;

		inst_bytes	[259][0]	= 8'hFF;
		inst_bytes	[259][1]	= 8'hC1;
		inst_size	[259]		= 4'd2;

		inst_bytes	[260][0]	= 8'hFF;
		inst_bytes	[260][1]	= 8'h01;
		inst_size	[260]		= 4'd2;

		inst_bytes	[261][0]	= 8'hFF;
		inst_bytes	[261][1]	= 8'h04;
		inst_bytes	[261][2]	= 8'h52;
		inst_size	[261]		= 4'd3;

		inst_bytes	[262][0]	= 8'hFF;
		inst_bytes	[262][1]	= 8'h05;
		inst_bytes	[262][2]	= 8'h01;
		inst_bytes	[262][3]	= 8'h02;
		inst_bytes	[262][4]	= 8'h03;
		inst_bytes	[262][5]	= 8'h04;
		inst_size	[262]		= 4'd6;

		inst_bytes	[263][0]	= 8'hFF;
		inst_bytes	[263][1]	= 8'h41;
		inst_bytes	[263][2]	= 8'h01;
		inst_size	[263]		= 4'd3;

		inst_bytes	[264][0]	= 8'hFF;
		inst_bytes	[264][1]	= 8'h44;
		inst_bytes	[264][2]	= 8'h52;
		inst_bytes	[264][3]	= 8'h01;
		inst_size	[264]		= 4'd4;

		inst_bytes	[265][0]	= 8'hFF;
		inst_bytes	[265][1]	= 8'h81;
		inst_bytes	[265][2]	= 8'h01;
		inst_bytes	[265][3]	= 8'h02;
		inst_bytes	[265][4]	= 8'h03;
		inst_bytes	[265][5]	= 8'h04;
		inst_size	[265]		= 4'd6;

		inst_bytes	[266][0]	= 8'hFF;
		inst_bytes	[266][1]	= 8'h84;
		inst_bytes	[266][2]	= 8'h52;
		inst_bytes	[266][3]	= 8'h01;
		inst_bytes	[266][4]	= 8'h02;
		inst_bytes	[266][5]	= 8'h03;
		inst_bytes	[266][6]	= 8'h04;
		inst_size	[266]		= 4'd7;

		inst_bytes	[267][0]	= 8'hFF;
		inst_bytes	[267][1]	= 8'hC1;
		inst_size	[267]		= 4'd2;

		inst_bytes	[268][0]	= 8'h66;
		inst_bytes	[268][1]	= 8'h41;
		inst_size	[268]		= 4'd2;

		inst_bytes	[269][0]	= 8'h41;
		inst_size	[269]		= 4'd1;

		inst_bytes	[270][0]	= 8'hCF;
		inst_size	[270]		= 4'd1;

		inst_bytes	[271][0]	= 8'h77;
		inst_bytes	[271][1]	= 8'h11;
		inst_size	[271]		= 4'd2;

		inst_bytes	[272][0]	= 8'h75;
		inst_bytes	[272][1]	= 8'h11;
		inst_size	[272]		= 4'd2;

		inst_bytes	[273][0]	= 8'h66;
		inst_bytes	[273][1]	= 8'h0F;
		inst_bytes	[273][2]	= 8'h87;
		inst_bytes	[273][3]	= 8'h11;
		inst_bytes	[273][4]	= 8'h12;
		inst_size	[273]		= 4'd5;

		inst_bytes	[274][0]	= 8'h0F;
		inst_bytes	[274][1]	= 8'h87;
		inst_bytes	[274][2]	= 8'h11;
		inst_bytes	[274][3]	= 8'h12;
		inst_bytes	[274][4]	= 8'h13;
		inst_bytes	[274][5]	= 8'h14;
		inst_size	[274]		= 4'd6;

		inst_bytes	[275][0]	= 8'h66;
		inst_bytes	[275][1]	= 8'h0F;
		inst_bytes	[275][2]	= 8'h85;
		inst_bytes	[275][3]	= 8'h11;
		inst_bytes	[275][4]	= 8'h12;
		inst_size	[275]		= 4'd5;

		inst_bytes	[276][0]	= 8'h0F;
		inst_bytes	[276][1]	= 8'h85;
		inst_bytes	[276][2]	= 8'h11;
		inst_bytes	[276][3]	= 8'h12;
		inst_bytes	[276][4]	= 8'h13;
		inst_bytes	[276][5]	= 8'h14;
		inst_size	[276]		= 4'd6;

		inst_bytes	[277][0]	= 8'hEB;
		inst_bytes	[277][1]	= 8'h11;
		inst_size	[277]		= 4'd2;

		inst_bytes	[278][0]	= 8'h66;
		inst_bytes	[278][1]	= 8'hE9;
		inst_bytes	[278][2]	= 8'h11;
		inst_bytes	[278][3]	= 8'h12;
		inst_size	[278]		= 4'd4;

		inst_bytes	[279][0]	= 8'hE9;
		inst_bytes	[279][1]	= 8'h11;
		inst_bytes	[279][2]	= 8'h12;
		inst_bytes	[279][3]	= 8'h13;
		inst_bytes	[279][4]	= 8'h14;
		inst_size	[279]		= 4'd5;

		inst_bytes	[280][0]	= 8'hFF;
		inst_bytes	[280][1]	= 8'h21;
		inst_size	[280]		= 4'd2;

		inst_bytes	[281][0]	= 8'hFF;
		inst_bytes	[281][1]	= 8'h24;
		inst_bytes	[281][2]	= 8'h52;
		inst_size	[281]		= 4'd3;

		inst_bytes	[282][0]	= 8'hFF;
		inst_bytes	[282][1]	= 8'h25;
		inst_bytes	[282][2]	= 8'h01;
		inst_bytes	[282][3]	= 8'h02;
		inst_bytes	[282][4]	= 8'h03;
		inst_bytes	[282][5]	= 8'h04;
		inst_size	[282]		= 4'd6;

		inst_bytes	[283][0]	= 8'hFF;
		inst_bytes	[283][1]	= 8'h61;
		inst_bytes	[283][2]	= 8'h01;
		inst_size	[283]		= 4'd3;

		inst_bytes	[284][0]	= 8'hFF;
		inst_bytes	[284][1]	= 8'h64;
		inst_bytes	[284][2]	= 8'h52;
		inst_bytes	[284][3]	= 8'h01;
		inst_size	[284]		= 4'd4;

		inst_bytes	[285][0]	= 8'hFF;
		inst_bytes	[285][1]	= 8'hA1;
		inst_bytes	[285][2]	= 8'h01;
		inst_bytes	[285][3]	= 8'h02;
		inst_bytes	[285][4]	= 8'h03;
		inst_bytes	[285][5]	= 8'h04;
		inst_size	[285]		= 4'd6;

		inst_bytes	[286][0]	= 8'hFF;
		inst_bytes	[286][1]	= 8'hA4;
		inst_bytes	[286][2]	= 8'h52;
		inst_bytes	[286][3]	= 8'h01;
		inst_bytes	[286][4]	= 8'h02;
		inst_bytes	[286][5]	= 8'h03;
		inst_bytes	[286][6]	= 8'h04;
		inst_size	[286]		= 4'd7;

		inst_bytes	[287][0]	= 8'hFF;
		inst_bytes	[287][1]	= 8'hE1;
		inst_size	[287]		= 4'd2;

		inst_bytes	[288][0]	= 8'hFF;
		inst_bytes	[288][1]	= 8'h21;
		inst_size	[288]		= 4'd2;

		inst_bytes	[289][0]	= 8'hFF;
		inst_bytes	[289][1]	= 8'h24;
		inst_bytes	[289][2]	= 8'h52;
		inst_size	[289]		= 4'd3;

		inst_bytes	[290][0]	= 8'hFF;
		inst_bytes	[290][1]	= 8'h25;
		inst_bytes	[290][2]	= 8'h01;
		inst_bytes	[290][3]	= 8'h02;
		inst_bytes	[290][4]	= 8'h03;
		inst_bytes	[290][5]	= 8'h04;
		inst_size	[290]		= 4'd6;

		inst_bytes	[291][0]	= 8'hFF;
		inst_bytes	[291][1]	= 8'h61;
		inst_bytes	[291][2]	= 8'h01;
		inst_size	[291]		= 4'd3;

		inst_bytes	[292][0]	= 8'hFF;
		inst_bytes	[292][1]	= 8'h64;
		inst_bytes	[292][2]	= 8'h52;
		inst_bytes	[292][3]	= 8'h01;
		inst_size	[292]		= 4'd4;

		inst_bytes	[293][0]	= 8'hFF;
		inst_bytes	[293][1]	= 8'hA1;
		inst_bytes	[293][2]	= 8'h01;
		inst_bytes	[293][3]	= 8'h02;
		inst_bytes	[293][4]	= 8'h03;
		inst_bytes	[293][5]	= 8'h04;
		inst_size	[293]		= 4'd6;

		inst_bytes	[294][0]	= 8'hFF;
		inst_bytes	[294][1]	= 8'hA4;
		inst_bytes	[294][2]	= 8'h52;
		inst_bytes	[294][3]	= 8'h01;
		inst_bytes	[294][4]	= 8'h02;
		inst_bytes	[294][5]	= 8'h03;
		inst_bytes	[294][6]	= 8'h04;
		inst_size	[294]		= 4'd7;

		inst_bytes	[295][0]	= 8'hFF;
		inst_bytes	[295][1]	= 8'hE1;
		inst_size	[295]		= 4'd2;

		inst_bytes	[296][0]	= 8'h66;
		inst_bytes	[296][1]	= 8'hEA;
		inst_bytes	[296][2]	= 8'h11;
		inst_bytes	[296][3]	= 8'h12;
		inst_bytes	[296][4]	= 8'h13;
		inst_bytes	[296][5]	= 8'h14;
		inst_size	[296]		= 4'd6;

		inst_bytes	[297][0]	= 8'hEA;
		inst_bytes	[297][1]	= 8'h0F;
		inst_bytes	[297][2]	= 8'h10;
		inst_bytes	[297][3]	= 8'h11;
		inst_bytes	[297][4]	= 8'h12;
		inst_bytes	[297][5]	= 8'h13;
		inst_bytes	[297][6]	= 8'h14;
		inst_size	[297]		= 4'd7;

		inst_bytes	[298][0]	= 8'h88;
		inst_bytes	[298][1]	= 8'h01;
		inst_size	[298]		= 4'd2;

		inst_bytes	[299][0]	= 8'h88;
		inst_bytes	[299][1]	= 8'h04;
		inst_bytes	[299][2]	= 8'h52;
		inst_size	[299]		= 4'd3;

		inst_bytes	[300][0]	= 8'h88;
		inst_bytes	[300][1]	= 8'h05;
		inst_bytes	[300][2]	= 8'h01;
		inst_bytes	[300][3]	= 8'h02;
		inst_bytes	[300][4]	= 8'h03;
		inst_bytes	[300][5]	= 8'h04;
		inst_size	[300]		= 4'd6;

		inst_bytes	[301][0]	= 8'h88;
		inst_bytes	[301][1]	= 8'h41;
		inst_bytes	[301][2]	= 8'h01;
		inst_size	[301]		= 4'd3;

		inst_bytes	[302][0]	= 8'h88;
		inst_bytes	[302][1]	= 8'h44;
		inst_bytes	[302][2]	= 8'h52;
		inst_bytes	[302][3]	= 8'h01;
		inst_size	[302]		= 4'd4;

		inst_bytes	[303][0]	= 8'h88;
		inst_bytes	[303][1]	= 8'h81;
		inst_bytes	[303][2]	= 8'h01;
		inst_bytes	[303][3]	= 8'h02;
		inst_bytes	[303][4]	= 8'h03;
		inst_bytes	[303][5]	= 8'h04;
		inst_size	[303]		= 4'd6;

		inst_bytes	[304][0]	= 8'h88;
		inst_bytes	[304][1]	= 8'h84;
		inst_bytes	[304][2]	= 8'h52;
		inst_bytes	[304][3]	= 8'h01;
		inst_bytes	[304][4]	= 8'h02;
		inst_bytes	[304][5]	= 8'h03;
		inst_bytes	[304][6]	= 8'h04;
		inst_size	[304]		= 4'd7;

		inst_bytes	[305][0]	= 8'h88;
		inst_bytes	[305][1]	= 8'hC1;
		inst_size	[305]		= 4'd2;

		inst_bytes	[306][0]	= 8'h89;
		inst_bytes	[306][1]	= 8'h01;
		inst_size	[306]		= 4'd2;

		inst_bytes	[307][0]	= 8'h89;
		inst_bytes	[307][1]	= 8'h04;
		inst_bytes	[307][2]	= 8'h52;
		inst_size	[307]		= 4'd3;

		inst_bytes	[308][0]	= 8'h89;
		inst_bytes	[308][1]	= 8'h05;
		inst_bytes	[308][2]	= 8'h01;
		inst_bytes	[308][3]	= 8'h02;
		inst_bytes	[308][4]	= 8'h03;
		inst_bytes	[308][5]	= 8'h04;
		inst_size	[308]		= 4'd6;

		inst_bytes	[309][0]	= 8'h89;
		inst_bytes	[309][1]	= 8'h41;
		inst_bytes	[309][2]	= 8'h01;
		inst_size	[309]		= 4'd3;

		inst_bytes	[310][0]	= 8'h89;
		inst_bytes	[310][1]	= 8'h44;
		inst_bytes	[310][2]	= 8'h52;
		inst_bytes	[310][3]	= 8'h01;
		inst_size	[310]		= 4'd4;

		inst_bytes	[311][0]	= 8'h89;
		inst_bytes	[311][1]	= 8'h81;
		inst_bytes	[311][2]	= 8'h01;
		inst_bytes	[311][3]	= 8'h02;
		inst_bytes	[311][4]	= 8'h03;
		inst_bytes	[311][5]	= 8'h04;
		inst_size	[311]		= 4'd6;

		inst_bytes	[312][0]	= 8'h89;
		inst_bytes	[312][1]	= 8'h84;
		inst_bytes	[312][2]	= 8'h52;
		inst_bytes	[312][3]	= 8'h01;
		inst_bytes	[312][4]	= 8'h02;
		inst_bytes	[312][5]	= 8'h03;
		inst_bytes	[312][6]	= 8'h04;
		inst_size	[312]		= 4'd7;

		inst_bytes	[313][0]	= 8'h89;
		inst_bytes	[313][1]	= 8'hC1;
		inst_size	[313]		= 4'd2;

		inst_bytes	[314][0]	= 8'h89;
		inst_bytes	[314][1]	= 8'h01;
		inst_size	[314]		= 4'd2;

		inst_bytes	[315][0]	= 8'h89;
		inst_bytes	[315][1]	= 8'h04;
		inst_bytes	[315][2]	= 8'h52;
		inst_size	[315]		= 4'd3;

		inst_bytes	[316][0]	= 8'h89;
		inst_bytes	[316][1]	= 8'h05;
		inst_bytes	[316][2]	= 8'h01;
		inst_bytes	[316][3]	= 8'h02;
		inst_bytes	[316][4]	= 8'h03;
		inst_bytes	[316][5]	= 8'h04;
		inst_size	[316]		= 4'd6;

		inst_bytes	[317][0]	= 8'h89;
		inst_bytes	[317][1]	= 8'h41;
		inst_bytes	[317][2]	= 8'h01;
		inst_size	[317]		= 4'd3;

		inst_bytes	[318][0]	= 8'h89;
		inst_bytes	[318][1]	= 8'h44;
		inst_bytes	[318][2]	= 8'h52;
		inst_bytes	[318][3]	= 8'h01;
		inst_size	[318]		= 4'd4;

		inst_bytes	[319][0]	= 8'h89;
		inst_bytes	[319][1]	= 8'h81;
		inst_bytes	[319][2]	= 8'h01;
		inst_bytes	[319][3]	= 8'h02;
		inst_bytes	[319][4]	= 8'h03;
		inst_bytes	[319][5]	= 8'h04;
		inst_size	[319]		= 4'd6;

		inst_bytes	[320][0]	= 8'h89;
		inst_bytes	[320][1]	= 8'h84;
		inst_bytes	[320][2]	= 8'h52;
		inst_bytes	[320][3]	= 8'h01;
		inst_bytes	[320][4]	= 8'h02;
		inst_bytes	[320][5]	= 8'h03;
		inst_bytes	[320][6]	= 8'h04;
		inst_size	[320]		= 4'd7;

		inst_bytes	[321][0]	= 8'h89;
		inst_bytes	[321][1]	= 8'hC1;
		inst_size	[321]		= 4'd2;

		inst_bytes	[322][0]	= 8'h8A;
		inst_bytes	[322][1]	= 8'h01;
		inst_size	[322]		= 4'd2;

		inst_bytes	[323][0]	= 8'h8A;
		inst_bytes	[323][1]	= 8'h04;
		inst_bytes	[323][2]	= 8'h52;
		inst_size	[323]		= 4'd3;

		inst_bytes	[324][0]	= 8'h8A;
		inst_bytes	[324][1]	= 8'h05;
		inst_bytes	[324][2]	= 8'h01;
		inst_bytes	[324][3]	= 8'h02;
		inst_bytes	[324][4]	= 8'h03;
		inst_bytes	[324][5]	= 8'h04;
		inst_size	[324]		= 4'd6;

		inst_bytes	[325][0]	= 8'h8A;
		inst_bytes	[325][1]	= 8'h41;
		inst_bytes	[325][2]	= 8'h01;
		inst_size	[325]		= 4'd3;

		inst_bytes	[326][0]	= 8'h8A;
		inst_bytes	[326][1]	= 8'h44;
		inst_bytes	[326][2]	= 8'h52;
		inst_bytes	[326][3]	= 8'h01;
		inst_size	[326]		= 4'd4;

		inst_bytes	[327][0]	= 8'h8A;
		inst_bytes	[327][1]	= 8'h81;
		inst_bytes	[327][2]	= 8'h01;
		inst_bytes	[327][3]	= 8'h02;
		inst_bytes	[327][4]	= 8'h03;
		inst_bytes	[327][5]	= 8'h04;
		inst_size	[327]		= 4'd6;

		inst_bytes	[328][0]	= 8'h8A;
		inst_bytes	[328][1]	= 8'h84;
		inst_bytes	[328][2]	= 8'h52;
		inst_bytes	[328][3]	= 8'h01;
		inst_bytes	[328][4]	= 8'h02;
		inst_bytes	[328][5]	= 8'h03;
		inst_bytes	[328][6]	= 8'h04;
		inst_size	[328]		= 4'd7;

		inst_bytes	[329][0]	= 8'h8A;
		inst_bytes	[329][1]	= 8'hC1;
		inst_size	[329]		= 4'd2;

		inst_bytes	[330][0]	= 8'h8B;
		inst_bytes	[330][1]	= 8'h01;
		inst_size	[330]		= 4'd2;

		inst_bytes	[331][0]	= 8'h8B;
		inst_bytes	[331][1]	= 8'h04;
		inst_bytes	[331][2]	= 8'h52;
		inst_size	[331]		= 4'd3;

		inst_bytes	[332][0]	= 8'h8B;
		inst_bytes	[332][1]	= 8'h05;
		inst_bytes	[332][2]	= 8'h01;
		inst_bytes	[332][3]	= 8'h02;
		inst_bytes	[332][4]	= 8'h03;
		inst_bytes	[332][5]	= 8'h04;
		inst_size	[332]		= 4'd6;

		inst_bytes	[333][0]	= 8'h8B;
		inst_bytes	[333][1]	= 8'h41;
		inst_bytes	[333][2]	= 8'h01;
		inst_size	[333]		= 4'd3;

		inst_bytes	[334][0]	= 8'h8B;
		inst_bytes	[334][1]	= 8'h44;
		inst_bytes	[334][2]	= 8'h52;
		inst_bytes	[334][3]	= 8'h01;
		inst_size	[334]		= 4'd4;

		inst_bytes	[335][0]	= 8'h8B;
		inst_bytes	[335][1]	= 8'h81;
		inst_bytes	[335][2]	= 8'h01;
		inst_bytes	[335][3]	= 8'h02;
		inst_bytes	[335][4]	= 8'h03;
		inst_bytes	[335][5]	= 8'h04;
		inst_size	[335]		= 4'd6;

		inst_bytes	[336][0]	= 8'h8B;
		inst_bytes	[336][1]	= 8'h84;
		inst_bytes	[336][2]	= 8'h52;
		inst_bytes	[336][3]	= 8'h01;
		inst_bytes	[336][4]	= 8'h02;
		inst_bytes	[336][5]	= 8'h03;
		inst_bytes	[336][6]	= 8'h04;
		inst_size	[336]		= 4'd7;

		inst_bytes	[337][0]	= 8'h8B;
		inst_bytes	[337][1]	= 8'hC1;
		inst_size	[337]		= 4'd2;

		inst_bytes	[338][0]	= 8'h8B;
		inst_bytes	[338][1]	= 8'h01;
		inst_size	[338]		= 4'd2;

		inst_bytes	[339][0]	= 8'h8B;
		inst_bytes	[339][1]	= 8'h04;
		inst_bytes	[339][2]	= 8'h52;
		inst_size	[339]		= 4'd3;

		inst_bytes	[340][0]	= 8'h8B;
		inst_bytes	[340][1]	= 8'h05;
		inst_bytes	[340][2]	= 8'h01;
		inst_bytes	[340][3]	= 8'h02;
		inst_bytes	[340][4]	= 8'h03;
		inst_bytes	[340][5]	= 8'h04;
		inst_size	[340]		= 4'd6;

		inst_bytes	[341][0]	= 8'h8B;
		inst_bytes	[341][1]	= 8'h41;
		inst_bytes	[341][2]	= 8'h01;
		inst_size	[341]		= 4'd3;

		inst_bytes	[342][0]	= 8'h8B;
		inst_bytes	[342][1]	= 8'h44;
		inst_bytes	[342][2]	= 8'h52;
		inst_bytes	[342][3]	= 8'h01;
		inst_size	[342]		= 4'd4;

		inst_bytes	[343][0]	= 8'h8B;
		inst_bytes	[343][1]	= 8'h81;
		inst_bytes	[343][2]	= 8'h01;
		inst_bytes	[343][3]	= 8'h02;
		inst_bytes	[343][4]	= 8'h03;
		inst_bytes	[343][5]	= 8'h04;
		inst_size	[343]		= 4'd6;

		inst_bytes	[344][0]	= 8'h8B;
		inst_bytes	[344][1]	= 8'h84;
		inst_bytes	[344][2]	= 8'h52;
		inst_bytes	[344][3]	= 8'h01;
		inst_bytes	[344][4]	= 8'h02;
		inst_bytes	[344][5]	= 8'h03;
		inst_bytes	[344][6]	= 8'h04;
		inst_size	[344]		= 4'd7;

		inst_bytes	[345][0]	= 8'h8B;
		inst_bytes	[345][1]	= 8'hC1;
		inst_size	[345]		= 4'd2;

		inst_bytes	[346][0]	= 8'h8C;
		inst_bytes	[346][1]	= 8'h01;
		inst_size	[346]		= 4'd2;

		inst_bytes	[347][0]	= 8'h8C;
		inst_bytes	[347][1]	= 8'h04;
		inst_bytes	[347][2]	= 8'h52;
		inst_size	[347]		= 4'd3;

		inst_bytes	[348][0]	= 8'h8C;
		inst_bytes	[348][1]	= 8'h05;
		inst_bytes	[348][2]	= 8'h01;
		inst_bytes	[348][3]	= 8'h02;
		inst_bytes	[348][4]	= 8'h03;
		inst_bytes	[348][5]	= 8'h04;
		inst_size	[348]		= 4'd6;

		inst_bytes	[349][0]	= 8'h8C;
		inst_bytes	[349][1]	= 8'h41;
		inst_bytes	[349][2]	= 8'h01;
		inst_size	[349]		= 4'd3;

		inst_bytes	[350][0]	= 8'h8C;
		inst_bytes	[350][1]	= 8'h44;
		inst_bytes	[350][2]	= 8'h52;
		inst_bytes	[350][3]	= 8'h01;
		inst_size	[350]		= 4'd4;

		inst_bytes	[351][0]	= 8'h8C;
		inst_bytes	[351][1]	= 8'h81;
		inst_bytes	[351][2]	= 8'h01;
		inst_bytes	[351][3]	= 8'h02;
		inst_bytes	[351][4]	= 8'h03;
		inst_bytes	[351][5]	= 8'h04;
		inst_size	[351]		= 4'd6;

		inst_bytes	[352][0]	= 8'h8C;
		inst_bytes	[352][1]	= 8'h84;
		inst_bytes	[352][2]	= 8'h52;
		inst_bytes	[352][3]	= 8'h01;
		inst_bytes	[352][4]	= 8'h02;
		inst_bytes	[352][5]	= 8'h03;
		inst_bytes	[352][6]	= 8'h04;
		inst_size	[352]		= 4'd7;

		inst_bytes	[353][0]	= 8'h8C;
		inst_bytes	[353][1]	= 8'hC1;
		inst_size	[353]		= 4'd2;

		inst_bytes	[354][0]	= 8'h8E;
		inst_bytes	[354][1]	= 8'h01;
		inst_size	[354]		= 4'd2;

		inst_bytes	[355][0]	= 8'h8E;
		inst_bytes	[355][1]	= 8'h04;
		inst_bytes	[355][2]	= 8'h52;
		inst_size	[355]		= 4'd3;

		inst_bytes	[356][0]	= 8'h8E;
		inst_bytes	[356][1]	= 8'h05;
		inst_bytes	[356][2]	= 8'h01;
		inst_bytes	[356][3]	= 8'h02;
		inst_bytes	[356][4]	= 8'h03;
		inst_bytes	[356][5]	= 8'h04;
		inst_size	[356]		= 4'd6;

		inst_bytes	[357][0]	= 8'h8E;
		inst_bytes	[357][1]	= 8'h41;
		inst_bytes	[357][2]	= 8'h01;
		inst_size	[357]		= 4'd3;

		inst_bytes	[358][0]	= 8'h8E;
		inst_bytes	[358][1]	= 8'h44;
		inst_bytes	[358][2]	= 8'h52;
		inst_bytes	[358][3]	= 8'h01;
		inst_size	[358]		= 4'd4;

		inst_bytes	[359][0]	= 8'h8E;
		inst_bytes	[359][1]	= 8'h81;
		inst_bytes	[359][2]	= 8'h01;
		inst_bytes	[359][3]	= 8'h02;
		inst_bytes	[359][4]	= 8'h03;
		inst_bytes	[359][5]	= 8'h04;
		inst_size	[359]		= 4'd6;

		inst_bytes	[360][0]	= 8'h8E;
		inst_bytes	[360][1]	= 8'h84;
		inst_bytes	[360][2]	= 8'h52;
		inst_bytes	[360][3]	= 8'h01;
		inst_bytes	[360][4]	= 8'h02;
		inst_bytes	[360][5]	= 8'h03;
		inst_bytes	[360][6]	= 8'h04;
		inst_size	[360]		= 4'd7;

		inst_bytes	[361][0]	= 8'h8E;
		inst_bytes	[361][1]	= 8'hC1;
		inst_size	[361]		= 4'd2;

		inst_bytes	[362][0]	= 8'hB1;
		inst_bytes	[362][1]	= 8'h11;
		inst_size	[362]		= 4'd2;

		inst_bytes	[363][0]	= 8'h66;
		inst_bytes	[363][1]	= 8'hB9;
		inst_bytes	[363][2]	= 8'h11;
		inst_bytes	[363][3]	= 8'h12;
		inst_size	[363]		= 4'd4;

		inst_bytes	[364][0]	= 8'hB9;
		inst_bytes	[364][1]	= 8'h11;
		inst_bytes	[364][2]	= 8'h12;
		inst_bytes	[364][3]	= 8'h13;
		inst_bytes	[364][4]	= 8'h14;
		inst_size	[364]		= 4'd5;

		inst_bytes	[365][0]	= 8'hC6;
		inst_bytes	[365][1]	= 8'h01;
		inst_bytes	[365][2]	= 8'h11;
		inst_size	[365]		= 4'd3;

		inst_bytes	[366][0]	= 8'hC6;
		inst_bytes	[366][1]	= 8'h04;
		inst_bytes	[366][2]	= 8'h52;
		inst_bytes	[366][3]	= 8'h11;
		inst_size	[366]		= 4'd4;

		inst_bytes	[367][0]	= 8'hC6;
		inst_bytes	[367][1]	= 8'h05;
		inst_bytes	[367][2]	= 8'h01;
		inst_bytes	[367][3]	= 8'h02;
		inst_bytes	[367][4]	= 8'h03;
		inst_bytes	[367][5]	= 8'h04;
		inst_bytes	[367][6]	= 8'h11;
		inst_size	[367]		= 4'd7;

		inst_bytes	[368][0]	= 8'hC6;
		inst_bytes	[368][1]	= 8'h41;
		inst_bytes	[368][2]	= 8'h01;
		inst_bytes	[368][3]	= 8'h11;
		inst_size	[368]		= 4'd4;

		inst_bytes	[369][0]	= 8'hC6;
		inst_bytes	[369][1]	= 8'h44;
		inst_bytes	[369][2]	= 8'h52;
		inst_bytes	[369][3]	= 8'h01;
		inst_bytes	[369][4]	= 8'h11;
		inst_size	[369]		= 4'd5;

		inst_bytes	[370][0]	= 8'hC6;
		inst_bytes	[370][1]	= 8'h81;
		inst_bytes	[370][2]	= 8'h01;
		inst_bytes	[370][3]	= 8'h02;
		inst_bytes	[370][4]	= 8'h03;
		inst_bytes	[370][5]	= 8'h04;
		inst_bytes	[370][6]	= 8'h11;
		inst_size	[370]		= 4'd7;

		inst_bytes	[371][0]	= 8'hC6;
		inst_bytes	[371][1]	= 8'h84;
		inst_bytes	[371][2]	= 8'h52;
		inst_bytes	[371][3]	= 8'h01;
		inst_bytes	[371][4]	= 8'h02;
		inst_bytes	[371][5]	= 8'h03;
		inst_bytes	[371][6]	= 8'h04;
		inst_bytes	[371][7]	= 8'h11;
		inst_size	[371]		= 4'd8;

		inst_bytes	[372][0]	= 8'hC6;
		inst_bytes	[372][1]	= 8'hC1;
		inst_bytes	[372][2]	= 8'h11;
		inst_size	[372]		= 4'd3;

		inst_bytes	[373][0]	= 8'h66;
		inst_bytes	[373][1]	= 8'hC7;
		inst_bytes	[373][2]	= 8'h01;
		inst_bytes	[373][3]	= 8'h11;
		inst_bytes	[373][4]	= 8'h12;
		inst_size	[373]		= 4'd5;

		inst_bytes	[374][0]	= 8'h66;
		inst_bytes	[374][1]	= 8'hC7;
		inst_bytes	[374][2]	= 8'h04;
		inst_bytes	[374][3]	= 8'h52;
		inst_bytes	[374][4]	= 8'h11;
		inst_bytes	[374][5]	= 8'h12;
		inst_size	[374]		= 4'd6;

		inst_bytes	[375][0]	= 8'h66;
		inst_bytes	[375][1]	= 8'hC7;
		inst_bytes	[375][2]	= 8'h05;
		inst_bytes	[375][3]	= 8'h01;
		inst_bytes	[375][4]	= 8'h02;
		inst_bytes	[375][5]	= 8'h03;
		inst_bytes	[375][6]	= 8'h04;
		inst_bytes	[375][7]	= 8'h11;
		inst_bytes	[375][8]	= 8'h12;
		inst_size	[375]		= 4'd9;

		inst_bytes	[376][0]	= 8'h66;
		inst_bytes	[376][1]	= 8'hC7;
		inst_bytes	[376][2]	= 8'h41;
		inst_bytes	[376][3]	= 8'h01;
		inst_bytes	[376][4]	= 8'h11;
		inst_bytes	[376][5]	= 8'h12;
		inst_size	[376]		= 4'd6;

		inst_bytes	[377][0]	= 8'h66;
		inst_bytes	[377][1]	= 8'hC7;
		inst_bytes	[377][2]	= 8'h44;
		inst_bytes	[377][3]	= 8'h52;
		inst_bytes	[377][4]	= 8'h01;
		inst_bytes	[377][5]	= 8'h11;
		inst_bytes	[377][6]	= 8'h12;
		inst_size	[377]		= 4'd7;

		inst_bytes	[378][0]	= 8'h66;
		inst_bytes	[378][1]	= 8'hC7;
		inst_bytes	[378][2]	= 8'h81;
		inst_bytes	[378][3]	= 8'h01;
		inst_bytes	[378][4]	= 8'h02;
		inst_bytes	[378][5]	= 8'h03;
		inst_bytes	[378][6]	= 8'h04;
		inst_bytes	[378][7]	= 8'h11;
		inst_bytes	[378][8]	= 8'h12;
		inst_size	[378]		= 4'd9;

		inst_bytes	[379][0]	= 8'h66;
		inst_bytes	[379][1]	= 8'hC7;
		inst_bytes	[379][2]	= 8'h84;
		inst_bytes	[379][3]	= 8'h52;
		inst_bytes	[379][4]	= 8'h01;
		inst_bytes	[379][5]	= 8'h02;
		inst_bytes	[379][6]	= 8'h03;
		inst_bytes	[379][7]	= 8'h04;
		inst_bytes	[379][8]	= 8'h11;
		inst_bytes	[379][9]	= 8'h12;
		inst_size	[379]		= 4'd10;

		inst_bytes	[380][0]	= 8'h66;
		inst_bytes	[380][1]	= 8'hC7;
		inst_bytes	[380][2]	= 8'hC1;
		inst_bytes	[380][3]	= 8'h11;
		inst_bytes	[380][4]	= 8'h12;
		inst_size	[380]		= 4'd5;

		inst_bytes	[381][0]	= 8'hC7;
		inst_bytes	[381][1]	= 8'h01;
		inst_bytes	[381][2]	= 8'h11;
		inst_bytes	[381][3]	= 8'h12;
		inst_bytes	[381][4]	= 8'h13;
		inst_bytes	[381][5]	= 8'h14;
		inst_size	[381]		= 4'd6;

		inst_bytes	[382][0]	= 8'hC7;
		inst_bytes	[382][1]	= 8'h04;
		inst_bytes	[382][2]	= 8'h52;
		inst_bytes	[382][3]	= 8'h11;
		inst_bytes	[382][4]	= 8'h12;
		inst_bytes	[382][5]	= 8'h13;
		inst_bytes	[382][6]	= 8'h14;
		inst_size	[382]		= 4'd7;

		inst_bytes	[383][0]	= 8'hC7;
		inst_bytes	[383][1]	= 8'h05;
		inst_bytes	[383][2]	= 8'h01;
		inst_bytes	[383][3]	= 8'h02;
		inst_bytes	[383][4]	= 8'h03;
		inst_bytes	[383][5]	= 8'h04;
		inst_bytes	[383][6]	= 8'h11;
		inst_bytes	[383][7]	= 8'h12;
		inst_bytes	[383][8]	= 8'h13;
		inst_bytes	[383][9]	= 8'h14;
		inst_size	[383]		= 4'd10;

		inst_bytes	[384][0]	= 8'hC7;
		inst_bytes	[384][1]	= 8'h41;
		inst_bytes	[384][2]	= 8'h01;
		inst_bytes	[384][3]	= 8'h11;
		inst_bytes	[384][4]	= 8'h12;
		inst_bytes	[384][5]	= 8'h13;
		inst_bytes	[384][6]	= 8'h14;
		inst_size	[384]		= 4'd7;

		inst_bytes	[385][0]	= 8'hC7;
		inst_bytes	[385][1]	= 8'h44;
		inst_bytes	[385][2]	= 8'h52;
		inst_bytes	[385][3]	= 8'h01;
		inst_bytes	[385][4]	= 8'h11;
		inst_bytes	[385][5]	= 8'h12;
		inst_bytes	[385][6]	= 8'h13;
		inst_bytes	[385][7]	= 8'h14;
		inst_size	[385]		= 4'd8;

		inst_bytes	[386][0]	= 8'hC7;
		inst_bytes	[386][1]	= 8'h81;
		inst_bytes	[386][2]	= 8'h01;
		inst_bytes	[386][3]	= 8'h02;
		inst_bytes	[386][4]	= 8'h03;
		inst_bytes	[386][5]	= 8'h04;
		inst_bytes	[386][6]	= 8'h11;
		inst_bytes	[386][7]	= 8'h12;
		inst_bytes	[386][8]	= 8'h13;
		inst_bytes	[386][9]	= 8'h14;
		inst_size	[386]		= 4'd10;

		inst_bytes	[387][0]	= 8'hC7;
		inst_bytes	[387][1]	= 8'h84;
		inst_bytes	[387][2]	= 8'h52;
		inst_bytes	[387][3]	= 8'h01;
		inst_bytes	[387][4]	= 8'h02;
		inst_bytes	[387][5]	= 8'h03;
		inst_bytes	[387][6]	= 8'h04;
		inst_bytes	[387][7]	= 8'h11;
		inst_bytes	[387][8]	= 8'h12;
		inst_bytes	[387][9]	= 8'h13;
		inst_bytes	[387][10]	= 8'h14;
		inst_size	[387]		= 4'd11;

		inst_bytes	[388][0]	= 8'hC7;
		inst_bytes	[388][1]	= 8'hC1;
		inst_bytes	[388][2]	= 8'h11;
		inst_bytes	[388][3]	= 8'h12;
		inst_bytes	[388][4]	= 8'h13;
		inst_bytes	[388][5]	= 8'h14;
		inst_size	[388]		= 4'd6;

		inst_bytes	[389][0]	= 8'h0F;
		inst_bytes	[389][1]	= 8'h6F;
		inst_bytes	[389][2]	= 8'h01;
		inst_size	[389]		= 4'd3;

		inst_bytes	[390][0]	= 8'h0F;
		inst_bytes	[390][1]	= 8'h6F;
		inst_bytes	[390][2]	= 8'h04;
		inst_bytes	[390][3]	= 8'h52;
		inst_size	[390]		= 4'd4;

		inst_bytes	[391][0]	= 8'h0F;
		inst_bytes	[391][1]	= 8'h6F;
		inst_bytes	[391][2]	= 8'h05;
		inst_bytes	[391][3]	= 8'h01;
		inst_bytes	[391][4]	= 8'h02;
		inst_bytes	[391][5]	= 8'h03;
		inst_bytes	[391][6]	= 8'h04;
		inst_size	[391]		= 4'd7;

		inst_bytes	[392][0]	= 8'h0F;
		inst_bytes	[392][1]	= 8'h6F;
		inst_bytes	[392][2]	= 8'h41;
		inst_bytes	[392][3]	= 8'h01;
		inst_size	[392]		= 4'd4;

		inst_bytes	[393][0]	= 8'h0F;
		inst_bytes	[393][1]	= 8'h6F;
		inst_bytes	[393][2]	= 8'h44;
		inst_bytes	[393][3]	= 8'h52;
		inst_bytes	[393][4]	= 8'h01;
		inst_size	[393]		= 4'd5;

		inst_bytes	[394][0]	= 8'h0F;
		inst_bytes	[394][1]	= 8'h6F;
		inst_bytes	[394][2]	= 8'h81;
		inst_bytes	[394][3]	= 8'h01;
		inst_bytes	[394][4]	= 8'h02;
		inst_bytes	[394][5]	= 8'h03;
		inst_bytes	[394][6]	= 8'h04;
		inst_size	[394]		= 4'd7;

		inst_bytes	[395][0]	= 8'h0F;
		inst_bytes	[395][1]	= 8'h6F;
		inst_bytes	[395][2]	= 8'h84;
		inst_bytes	[395][3]	= 8'h52;
		inst_bytes	[395][4]	= 8'h01;
		inst_bytes	[395][5]	= 8'h02;
		inst_bytes	[395][6]	= 8'h03;
		inst_bytes	[395][7]	= 8'h04;
		inst_size	[395]		= 4'd8;

		inst_bytes	[396][0]	= 8'h0F;
		inst_bytes	[396][1]	= 8'h6F;
		inst_bytes	[396][2]	= 8'hC1;
		inst_size	[396]		= 4'd3;

		inst_bytes	[397][0]	= 8'h0F;
		inst_bytes	[397][1]	= 8'h7F;
		inst_bytes	[397][2]	= 8'h01;
		inst_size	[397]		= 4'd3;

		inst_bytes	[398][0]	= 8'h0F;
		inst_bytes	[398][1]	= 8'h7F;
		inst_bytes	[398][2]	= 8'h04;
		inst_bytes	[398][3]	= 8'h52;
		inst_size	[398]		= 4'd4;

		inst_bytes	[399][0]	= 8'h0F;
		inst_bytes	[399][1]	= 8'h7F;
		inst_bytes	[399][2]	= 8'h05;
		inst_bytes	[399][3]	= 8'h01;
		inst_bytes	[399][4]	= 8'h02;
		inst_bytes	[399][5]	= 8'h03;
		inst_bytes	[399][6]	= 8'h04;
		inst_size	[399]		= 4'd7;

		inst_bytes	[400][0]	= 8'h0F;
		inst_bytes	[400][1]	= 8'h7F;
		inst_bytes	[400][2]	= 8'h41;
		inst_bytes	[400][3]	= 8'h01;
		inst_size	[400]		= 4'd4;

		inst_bytes	[401][0]	= 8'h0F;
		inst_bytes	[401][1]	= 8'h7F;
		inst_bytes	[401][2]	= 8'h44;
		inst_bytes	[401][3]	= 8'h52;
		inst_bytes	[401][4]	= 8'h01;
		inst_size	[401]		= 4'd5;

		inst_bytes	[402][0]	= 8'h0F;
		inst_bytes	[402][1]	= 8'h7F;
		inst_bytes	[402][2]	= 8'h81;
		inst_bytes	[402][3]	= 8'h01;
		inst_bytes	[402][4]	= 8'h02;
		inst_bytes	[402][5]	= 8'h03;
		inst_bytes	[402][6]	= 8'h04;
		inst_size	[402]		= 4'd7;

		inst_bytes	[403][0]	= 8'h0F;
		inst_bytes	[403][1]	= 8'h7F;
		inst_bytes	[403][2]	= 8'h84;
		inst_bytes	[403][3]	= 8'h52;
		inst_bytes	[403][4]	= 8'h01;
		inst_bytes	[403][5]	= 8'h02;
		inst_bytes	[403][6]	= 8'h03;
		inst_bytes	[403][7]	= 8'h04;
		inst_size	[403]		= 4'd8;

		inst_bytes	[404][0]	= 8'h0F;
		inst_bytes	[404][1]	= 8'h7F;
		inst_bytes	[404][2]	= 8'hC1;
		inst_size	[404]		= 4'd3;

		inst_bytes	[405][0]	= 8'hF6;
		inst_bytes	[405][1]	= 8'h11;
		inst_size	[405]		= 4'd2;

		inst_bytes	[406][0]	= 8'hF6;
		inst_bytes	[406][1]	= 8'h14;
		inst_bytes	[406][2]	= 8'h52;
		inst_size	[406]		= 4'd3;

		inst_bytes	[407][0]	= 8'hF6;
		inst_bytes	[407][1]	= 8'h15;
		inst_bytes	[407][2]	= 8'h01;
		inst_bytes	[407][3]	= 8'h02;
		inst_bytes	[407][4]	= 8'h03;
		inst_bytes	[407][5]	= 8'h04;
		inst_size	[407]		= 4'd6;

		inst_bytes	[408][0]	= 8'hF6;
		inst_bytes	[408][1]	= 8'h51;
		inst_bytes	[408][2]	= 8'h01;
		inst_size	[408]		= 4'd3;

		inst_bytes	[409][0]	= 8'hF6;
		inst_bytes	[409][1]	= 8'h54;
		inst_bytes	[409][2]	= 8'h52;
		inst_bytes	[409][3]	= 8'h01;
		inst_size	[409]		= 4'd4;

		inst_bytes	[410][0]	= 8'hF6;
		inst_bytes	[410][1]	= 8'h91;
		inst_bytes	[410][2]	= 8'h01;
		inst_bytes	[410][3]	= 8'h02;
		inst_bytes	[410][4]	= 8'h04;
		inst_bytes	[410][5]	= 8'h04;
		inst_size	[410]		= 4'd6;

		inst_bytes	[411][0]	= 8'hF6;
		inst_bytes	[411][1]	= 8'h94;
		inst_bytes	[411][2]	= 8'h52;
		inst_bytes	[411][3]	= 8'h01;
		inst_bytes	[411][4]	= 8'h02;
		inst_bytes	[411][5]	= 8'h03;
		inst_bytes	[411][6]	= 8'h04;
		inst_size	[411]		= 4'd7;

		inst_bytes	[412][0]	= 8'hF6;
		inst_bytes	[412][1]	= 8'hD1;
		inst_size	[412]		= 4'd2;

		inst_bytes	[413][0]	= 8'hF7;
		inst_bytes	[413][1]	= 8'h11;
		inst_size	[413]		= 4'd2;

		inst_bytes	[414][0]	= 8'hF7;
		inst_bytes	[414][1]	= 8'h14;
		inst_bytes	[414][2]	= 8'h52;
		inst_size	[414]		= 4'd3;

		inst_bytes	[415][0]	= 8'hF7;
		inst_bytes	[415][1]	= 8'h15;
		inst_bytes	[415][2]	= 8'h01;
		inst_bytes	[415][3]	= 8'h02;
		inst_bytes	[415][4]	= 8'h03;
		inst_bytes	[415][5]	= 8'h04;
		inst_size	[415]		= 4'd6;

		inst_bytes	[416][0]	= 8'hF7;
		inst_bytes	[416][1]	= 8'h51;
		inst_bytes	[416][2]	= 8'h01;
		inst_size	[416]		= 4'd3;

		inst_bytes	[417][0]	= 8'hF7;
		inst_bytes	[417][1]	= 8'h54;
		inst_bytes	[417][2]	= 8'h52;
		inst_bytes	[417][3]	= 8'h01;
		inst_size	[417]		= 4'd4;

		inst_bytes	[418][0]	= 8'hF7;
		inst_bytes	[418][1]	= 8'h91;
		inst_bytes	[418][2]	= 8'h01;
		inst_bytes	[418][3]	= 8'h02;
		inst_bytes	[418][4]	= 8'h04;
		inst_bytes	[418][5]	= 8'h04;
		inst_size	[418]		= 4'd6;

		inst_bytes	[419][0]	= 8'hF7;
		inst_bytes	[419][1]	= 8'h94;
		inst_bytes	[419][2]	= 8'h52;
		inst_bytes	[419][3]	= 8'h01;
		inst_bytes	[419][4]	= 8'h02;
		inst_bytes	[419][5]	= 8'h03;
		inst_bytes	[419][6]	= 8'h04;
		inst_size	[419]		= 4'd7;

		inst_bytes	[420][0]	= 8'hF7;
		inst_bytes	[420][1]	= 8'hD1;
		inst_size	[420]		= 4'd2;

		inst_bytes	[421][0]	= 8'hF7;
		inst_bytes	[421][1]	= 8'h11;
		inst_size	[421]		= 4'd2;

		inst_bytes	[422][0]	= 8'hF7;
		inst_bytes	[422][1]	= 8'h14;
		inst_bytes	[422][2]	= 8'h52;
		inst_size	[422]		= 4'd3;

		inst_bytes	[423][0]	= 8'hF7;
		inst_bytes	[423][1]	= 8'h15;
		inst_bytes	[423][2]	= 8'h01;
		inst_bytes	[423][3]	= 8'h02;
		inst_bytes	[423][4]	= 8'h03;
		inst_bytes	[423][5]	= 8'h04;
		inst_size	[423]		= 4'd6;

		inst_bytes	[424][0]	= 8'hF7;
		inst_bytes	[424][1]	= 8'h51;
		inst_bytes	[424][2]	= 8'h01;
		inst_size	[424]		= 4'd3;

		inst_bytes	[425][0]	= 8'hF7;
		inst_bytes	[425][1]	= 8'h54;
		inst_bytes	[425][2]	= 8'h52;
		inst_bytes	[425][3]	= 8'h01;
		inst_size	[425]		= 4'd4;

		inst_bytes	[426][0]	= 8'hF7;
		inst_bytes	[426][1]	= 8'h91;
		inst_bytes	[426][2]	= 8'h01;
		inst_bytes	[426][3]	= 8'h02;
		inst_bytes	[426][4]	= 8'h04;
		inst_bytes	[426][5]	= 8'h04;
		inst_size	[426]		= 4'd6;

		inst_bytes	[427][0]	= 8'hF7;
		inst_bytes	[427][1]	= 8'h94;
		inst_bytes	[427][2]	= 8'h52;
		inst_bytes	[427][3]	= 8'h01;
		inst_bytes	[427][4]	= 8'h02;
		inst_bytes	[427][5]	= 8'h03;
		inst_bytes	[427][6]	= 8'h04;
		inst_size	[427]		= 4'd7;

		inst_bytes	[428][0]	= 8'hF7;
		inst_bytes	[428][1]	= 8'hD1;
		inst_size	[428]		= 4'd2;

		inst_bytes	[429][0]	= 8'h0C;
		inst_bytes	[429][1]	= 8'h11;
		inst_size	[429]		= 4'd2;

		inst_bytes	[430][0]	= 8'h66;
		inst_bytes	[430][1]	= 8'h0D;
		inst_bytes	[430][2]	= 8'h11;
		inst_bytes	[430][3]	= 8'h12;
		inst_size	[430]		= 4'd4;

		inst_bytes	[431][0]	= 8'h0D;
		inst_bytes	[431][1]	= 8'h11;
		inst_bytes	[431][2]	= 8'h12;
		inst_bytes	[431][3]	= 8'h13;
		inst_bytes	[431][4]	= 8'h14;
		inst_size	[431]		= 4'd5;

		inst_bytes	[432][0]	= 8'h80;
		inst_bytes	[432][1]	= 8'h09;
		inst_bytes	[432][2]	= 8'h11;
		inst_size	[432]		= 4'd3;

		inst_bytes	[433][0]	= 8'h80;
		inst_bytes	[433][1]	= 8'h0C;
		inst_bytes	[433][2]	= 8'h52;
		inst_bytes	[433][3]	= 8'h11;
		inst_size	[433]		= 4'd4;

		inst_bytes	[434][0]	= 8'h80;
		inst_bytes	[434][1]	= 8'h0D;
		inst_bytes	[434][2]	= 8'h01;
		inst_bytes	[434][3]	= 8'h02;
		inst_bytes	[434][4]	= 8'h03;
		inst_bytes	[434][5]	= 8'h04;
		inst_bytes	[434][6]	= 8'h11;
		inst_size	[434]		= 4'd7;

		inst_bytes	[435][0]	= 8'h80;
		inst_bytes	[435][1]	= 8'h49;
		inst_bytes	[435][2]	= 8'h01;
		inst_bytes	[435][3]	= 8'h11;
		inst_size	[435]		= 4'd4;

		inst_bytes	[436][0]	= 8'h80;
		inst_bytes	[436][1]	= 8'h4C;
		inst_bytes	[436][2]	= 8'h52;
		inst_bytes	[436][3]	= 8'h01;
		inst_bytes	[436][4]	= 8'h11;
		inst_size	[436]		= 4'd5;

		inst_bytes	[437][0]	= 8'h80;
		inst_bytes	[437][1]	= 8'h89;
		inst_bytes	[437][2]	= 8'h01;
		inst_bytes	[437][3]	= 8'h02;
		inst_bytes	[437][4]	= 8'h03;
		inst_bytes	[437][5]	= 8'h04;
		inst_bytes	[437][6]	= 8'h11;
		inst_size	[437]		= 4'd7;

		inst_bytes	[438][0]	= 8'h80;
		inst_bytes	[438][1]	= 8'h8C;
		inst_bytes	[438][2]	= 8'h52;
		inst_bytes	[438][3]	= 8'h01;
		inst_bytes	[438][4]	= 8'h02;
		inst_bytes	[438][5]	= 8'h03;
		inst_bytes	[438][6]	= 8'h04;
		inst_bytes	[438][7]	= 8'h11;
		inst_size	[438]		= 4'd8;

		inst_bytes	[439][0]	= 8'h80;
		inst_bytes	[439][1]	= 8'hC9;
		inst_bytes	[439][2]	= 8'h11;
		inst_size	[439]		= 4'd3;

		inst_bytes	[440][0]	= 8'h66;
		inst_bytes	[440][1]	= 8'h81;
		inst_bytes	[440][2]	= 8'h09;
		inst_bytes	[440][3]	= 8'h11;
		inst_bytes	[440][4]	= 8'h12;
		inst_size	[440]		= 4'd5;

		inst_bytes	[441][0]	= 8'h66;
		inst_bytes	[441][1]	= 8'h81;
		inst_bytes	[441][2]	= 8'h0C;
		inst_bytes	[441][3]	= 8'h52;
		inst_bytes	[441][4]	= 8'h11;
		inst_bytes	[441][5]	= 8'h12;
		inst_size	[441]		= 4'd6;

		inst_bytes	[442][0]	= 8'h66;
		inst_bytes	[442][1]	= 8'h81;
		inst_bytes	[442][2]	= 8'h0D;
		inst_bytes	[442][3]	= 8'h01;
		inst_bytes	[442][4]	= 8'h02;
		inst_bytes	[442][5]	= 8'h03;
		inst_bytes	[442][6]	= 8'h04;
		inst_bytes	[442][7]	= 8'h11;
		inst_bytes	[442][8]	= 8'h12;
		inst_size	[442]		= 4'd9;

		inst_bytes	[443][0]	= 8'h66;
		inst_bytes	[443][1]	= 8'h81;
		inst_bytes	[443][2]	= 8'h49;
		inst_bytes	[443][3]	= 8'h01;
		inst_bytes	[443][4]	= 8'h11;
		inst_bytes	[443][5]	= 8'h12;
		inst_size	[443]		= 4'd6;

		inst_bytes	[444][0]	= 8'h66;
		inst_bytes	[444][1]	= 8'h81;
		inst_bytes	[444][2]	= 8'h4C;
		inst_bytes	[444][3]	= 8'h52;
		inst_bytes	[444][4]	= 8'h01;
		inst_bytes	[444][5]	= 8'h11;
		inst_bytes	[444][6]	= 8'h12;
		inst_size	[444]		= 4'd7;

		inst_bytes	[445][0]	= 8'h66;
		inst_bytes	[445][1]	= 8'h81;
		inst_bytes	[445][2]	= 8'h89;
		inst_bytes	[445][3]	= 8'h01;
		inst_bytes	[445][4]	= 8'h02;
		inst_bytes	[445][5]	= 8'h03;
		inst_bytes	[445][6]	= 8'h04;
		inst_bytes	[445][7]	= 8'h11;
		inst_bytes	[445][8]	= 8'h12;
		inst_size	[445]		= 4'd9;

		inst_bytes	[446][0]	= 8'h66;
		inst_bytes	[446][1]	= 8'h81;
		inst_bytes	[446][2]	= 8'h8C;
		inst_bytes	[446][3]	= 8'h52;
		inst_bytes	[446][4]	= 8'h01;
		inst_bytes	[446][5]	= 8'h02;
		inst_bytes	[446][6]	= 8'h03;
		inst_bytes	[446][7]	= 8'h04;
		inst_bytes	[446][8]	= 8'h11;
		inst_bytes	[446][9]	= 8'h12;
		inst_size	[446]		= 4'd10;

		inst_bytes	[447][0]	= 8'h66;
		inst_bytes	[447][1]	= 8'h81;
		inst_bytes	[447][2]	= 8'hC9;
		inst_bytes	[447][3]	= 8'h11;
		inst_bytes	[447][4]	= 8'h12;
		inst_size	[447]		= 4'd5;

		inst_bytes	[448][0]	= 8'h81;
		inst_bytes	[448][1]	= 8'h09;
		inst_bytes	[448][2]	= 8'h11;
		inst_bytes	[448][3]	= 8'h12;
		inst_bytes	[448][4]	= 8'h13;
		inst_bytes	[448][5]	= 8'h14;
		inst_size	[448]		= 4'd6;

		inst_bytes	[449][0]	= 8'h81;
		inst_bytes	[449][1]	= 8'h0C;
		inst_bytes	[449][2]	= 8'h52;
		inst_bytes	[449][3]	= 8'h11;
		inst_bytes	[449][4]	= 8'h12;
		inst_bytes	[449][5]	= 8'h13;
		inst_bytes	[449][6]	= 8'h14;
		inst_size	[449]		= 4'd7;

		inst_bytes	[450][0]	= 8'h81;
		inst_bytes	[450][1]	= 8'h0D;
		inst_bytes	[450][2]	= 8'h01;
		inst_bytes	[450][3]	= 8'h02;
		inst_bytes	[450][4]	= 8'h03;
		inst_bytes	[450][5]	= 8'h04;
		inst_bytes	[450][6]	= 8'h11;
		inst_bytes	[450][7]	= 8'h12;
		inst_bytes	[450][8]	= 8'h13;
		inst_bytes	[450][9]	= 8'h14;
		inst_size	[450]		= 4'd10;

		inst_bytes	[451][0]	= 8'h81;
		inst_bytes	[451][1]	= 8'h49;
		inst_bytes	[451][2]	= 8'h01;
		inst_bytes	[451][3]	= 8'h11;
		inst_bytes	[451][4]	= 8'h12;
		inst_bytes	[451][5]	= 8'h13;
		inst_bytes	[451][6]	= 8'h14;
		inst_size	[451]		= 4'd7;

		inst_bytes	[452][0]	= 8'h81;
		inst_bytes	[452][1]	= 8'h4C;
		inst_bytes	[452][2]	= 8'h52;
		inst_bytes	[452][3]	= 8'h01;
		inst_bytes	[452][4]	= 8'h11;
		inst_bytes	[452][5]	= 8'h12;
		inst_bytes	[452][6]	= 8'h13;
		inst_bytes	[452][7]	= 8'h14;
		inst_size	[452]		= 4'd8;

		inst_bytes	[453][0]	= 8'h81;
		inst_bytes	[453][1]	= 8'h89;
		inst_bytes	[453][2]	= 8'h01;
		inst_bytes	[453][3]	= 8'h02;
		inst_bytes	[453][4]	= 8'h03;
		inst_bytes	[453][5]	= 8'h04;
		inst_bytes	[453][6]	= 8'h11;
		inst_bytes	[453][7]	= 8'h12;
		inst_bytes	[453][8]	= 8'h13;
		inst_bytes	[453][9]	= 8'h14;
		inst_size	[453]		= 4'd10;

		inst_bytes	[454][0]	= 8'h81;
		inst_bytes	[454][1]	= 8'h8C;
		inst_bytes	[454][2]	= 8'h52;
		inst_bytes	[454][3]	= 8'h01;
		inst_bytes	[454][4]	= 8'h02;
		inst_bytes	[454][5]	= 8'h03;
		inst_bytes	[454][6]	= 8'h04;
		inst_bytes	[454][7]	= 8'h11;
		inst_bytes	[454][8]	= 8'h12;
		inst_bytes	[454][9]	= 8'h13;
		inst_bytes	[454][10]	= 8'h14;
		inst_size	[454]		= 4'd11;

		inst_bytes	[455][0]	= 8'h81;
		inst_bytes	[455][1]	= 8'hC9;
		inst_bytes	[455][2]	= 8'h11;
		inst_bytes	[455][3]	= 8'h12;
		inst_bytes	[455][4]	= 8'h13;
		inst_bytes	[455][5]	= 8'h14;
		inst_size	[455]		= 4'd6;

		inst_bytes	[456][0]	= 8'h83;
		inst_bytes	[456][1]	= 8'h09;
		inst_bytes	[456][2]	= 8'h11;
		inst_size	[456]		= 4'd3;

		inst_bytes	[457][0]	= 8'h83;
		inst_bytes	[457][1]	= 8'h0C;
		inst_bytes	[457][2]	= 8'h52;
		inst_bytes	[457][3]	= 8'h11;
		inst_size	[457]		= 4'd4;

		inst_bytes	[458][0]	= 8'h83;
		inst_bytes	[458][1]	= 8'h0D;
		inst_bytes	[458][2]	= 8'h01;
		inst_bytes	[458][3]	= 8'h02;
		inst_bytes	[458][4]	= 8'h03;
		inst_bytes	[458][5]	= 8'h04;
		inst_bytes	[458][6]	= 8'h11;
		inst_size	[458]		= 4'd7;

		inst_bytes	[459][0]	= 8'h83;
		inst_bytes	[459][1]	= 8'h49;
		inst_bytes	[459][2]	= 8'h01;
		inst_bytes	[459][3]	= 8'h11;
		inst_size	[459]		= 4'd4;

		inst_bytes	[460][0]	= 8'h83;
		inst_bytes	[460][1]	= 8'h4C;
		inst_bytes	[460][2]	= 8'h52;
		inst_bytes	[460][3]	= 8'h01;
		inst_bytes	[460][4]	= 8'h11;
		inst_size	[460]		= 4'd5;

		inst_bytes	[461][0]	= 8'h83;
		inst_bytes	[461][1]	= 8'h89;
		inst_bytes	[461][2]	= 8'h01;
		inst_bytes	[461][3]	= 8'h02;
		inst_bytes	[461][4]	= 8'h03;
		inst_bytes	[461][5]	= 8'h04;
		inst_bytes	[461][6]	= 8'h11;
		inst_size	[461]		= 4'd7;

		inst_bytes	[462][0]	= 8'h83;
		inst_bytes	[462][1]	= 8'h8C;
		inst_bytes	[462][2]	= 8'h52;
		inst_bytes	[462][3]	= 8'h01;
		inst_bytes	[462][4]	= 8'h02;
		inst_bytes	[462][5]	= 8'h03;
		inst_bytes	[462][6]	= 8'h04;
		inst_bytes	[462][7]	= 8'h11;
		inst_size	[462]		= 4'd8;

		inst_bytes	[463][0]	= 8'h83;
		inst_bytes	[463][1]	= 8'hC9;
		inst_bytes	[463][2]	= 8'h11;
		inst_size	[463]		= 4'd3;

		inst_bytes	[464][0]	= 8'h83;
		inst_bytes	[464][1]	= 8'h09;
		inst_bytes	[464][2]	= 8'h11;
		inst_size	[464]		= 4'd3;

		inst_bytes	[465][0]	= 8'h83;
		inst_bytes	[465][1]	= 8'h0C;
		inst_bytes	[465][2]	= 8'h52;
		inst_bytes	[465][3]	= 8'h11;
		inst_size	[465]		= 4'd4;

		inst_bytes	[466][0]	= 8'h83;
		inst_bytes	[466][1]	= 8'h0D;
		inst_bytes	[466][2]	= 8'h01;
		inst_bytes	[466][3]	= 8'h02;
		inst_bytes	[466][4]	= 8'h03;
		inst_bytes	[466][5]	= 8'h04;
		inst_bytes	[466][6]	= 8'h11;
		inst_size	[466]		= 4'd7;

		inst_bytes	[467][0]	= 8'h83;
		inst_bytes	[467][1]	= 8'h49;
		inst_bytes	[467][2]	= 8'h01;
		inst_bytes	[467][3]	= 8'h11;
		inst_size	[467]		= 4'd4;

		inst_bytes	[468][0]	= 8'h83;
		inst_bytes	[468][1]	= 8'h4C;
		inst_bytes	[468][2]	= 8'h52;
		inst_bytes	[468][3]	= 8'h01;
		inst_bytes	[468][4]	= 8'h11;
		inst_size	[468]		= 4'd5;

		inst_bytes	[469][0]	= 8'h83;
		inst_bytes	[469][1]	= 8'h89;
		inst_bytes	[469][2]	= 8'h01;
		inst_bytes	[469][3]	= 8'h02;
		inst_bytes	[469][4]	= 8'h03;
		inst_bytes	[469][5]	= 8'h04;
		inst_bytes	[469][6]	= 8'h11;
		inst_size	[469]		= 4'd7;

		inst_bytes	[470][0]	= 8'h83;
		inst_bytes	[470][1]	= 8'h8C;
		inst_bytes	[470][2]	= 8'h52;
		inst_bytes	[470][3]	= 8'h01;
		inst_bytes	[470][4]	= 8'h02;
		inst_bytes	[470][5]	= 8'h03;
		inst_bytes	[470][6]	= 8'h04;
		inst_bytes	[470][7]	= 8'h11;
		inst_size	[470]		= 4'd8;

		inst_bytes	[471][0]	= 8'h83;
		inst_bytes	[471][1]	= 8'hC9;
		inst_bytes	[471][2]	= 8'h11;
		inst_size	[471]		= 4'd3;

		inst_bytes	[472][0]	= 8'h08;
		inst_bytes	[472][1]	= 8'h01;
		inst_size	[472]		= 4'd2;

		inst_bytes	[473][0]	= 8'h08;
		inst_bytes	[473][1]	= 8'h04;
		inst_bytes	[473][2]	= 8'h52;
		inst_size	[473]		= 4'd3;

		inst_bytes	[474][0]	= 8'h08;
		inst_bytes	[474][1]	= 8'h05;
		inst_bytes	[474][2]	= 8'h01;
		inst_bytes	[474][3]	= 8'h02;
		inst_bytes	[474][4]	= 8'h03;
		inst_bytes	[474][5]	= 8'h04;
		inst_size	[474]		= 4'd6;

		inst_bytes	[475][0]	= 8'h08;
		inst_bytes	[475][1]	= 8'h41;
		inst_bytes	[475][2]	= 8'h01;
		inst_size	[475]		= 4'd3;

		inst_bytes	[476][0]	= 8'h08;
		inst_bytes	[476][1]	= 8'h44;
		inst_bytes	[476][2]	= 8'h52;
		inst_bytes	[476][3]	= 8'h01;
		inst_size	[476]		= 4'd4;

		inst_bytes	[477][0]	= 8'h08;
		inst_bytes	[477][1]	= 8'h81;
		inst_bytes	[477][2]	= 8'h01;
		inst_bytes	[477][3]	= 8'h02;
		inst_bytes	[477][4]	= 8'h03;
		inst_bytes	[477][5]	= 8'h04;
		inst_size	[477]		= 4'd6;

		inst_bytes	[478][0]	= 8'h08;
		inst_bytes	[478][1]	= 8'h84;
		inst_bytes	[478][2]	= 8'h52;
		inst_bytes	[478][3]	= 8'h01;
		inst_bytes	[478][4]	= 8'h02;
		inst_bytes	[478][5]	= 8'h03;
		inst_bytes	[478][6]	= 8'h04;
		inst_size	[478]		= 4'd7;

		inst_bytes	[479][0]	= 8'h08;
		inst_bytes	[479][1]	= 8'hC1;
		inst_size	[479]		= 4'd2;

		inst_bytes	[480][0]	= 8'h09;
		inst_bytes	[480][1]	= 8'h01;
		inst_size	[480]		= 4'd2;

		inst_bytes	[481][0]	= 8'h09;
		inst_bytes	[481][1]	= 8'h04;
		inst_bytes	[481][2]	= 8'h52;
		inst_size	[481]		= 4'd3;

		inst_bytes	[482][0]	= 8'h09;
		inst_bytes	[482][1]	= 8'h05;
		inst_bytes	[482][2]	= 8'h01;
		inst_bytes	[482][3]	= 8'h02;
		inst_bytes	[482][4]	= 8'h03;
		inst_bytes	[482][5]	= 8'h04;
		inst_size	[482]		= 4'd6;

		inst_bytes	[483][0]	= 8'h09;
		inst_bytes	[483][1]	= 8'h41;
		inst_bytes	[483][2]	= 8'h01;
		inst_size	[483]		= 4'd3;

		inst_bytes	[484][0]	= 8'h09;
		inst_bytes	[484][1]	= 8'h44;
		inst_bytes	[484][2]	= 8'h52;
		inst_bytes	[484][3]	= 8'h01;
		inst_size	[484]		= 4'd4;

		inst_bytes	[485][0]	= 8'h09;
		inst_bytes	[485][1]	= 8'h81;
		inst_bytes	[485][2]	= 8'h01;
		inst_bytes	[485][3]	= 8'h02;
		inst_bytes	[485][4]	= 8'h03;
		inst_bytes	[485][5]	= 8'h04;
		inst_size	[485]		= 4'd6;

		inst_bytes	[486][0]	= 8'h09;
		inst_bytes	[486][1]	= 8'h84;
		inst_bytes	[486][2]	= 8'h52;
		inst_bytes	[486][3]	= 8'h01;
		inst_bytes	[486][4]	= 8'h02;
		inst_bytes	[486][5]	= 8'h03;
		inst_bytes	[486][6]	= 8'h04;
		inst_size	[486]		= 4'd7;

		inst_bytes	[487][0]	= 8'h09;
		inst_bytes	[487][1]	= 8'hC1;
		inst_size	[487]		= 4'd2;

		inst_bytes	[488][0]	= 8'h09;
		inst_bytes	[488][1]	= 8'h01;
		inst_size	[488]		= 4'd2;

		inst_bytes	[489][0]	= 8'h09;
		inst_bytes	[489][1]	= 8'h04;
		inst_bytes	[489][2]	= 8'h52;
		inst_size	[489]		= 4'd3;

		inst_bytes	[490][0]	= 8'h09;
		inst_bytes	[490][1]	= 8'h05;
		inst_bytes	[490][2]	= 8'h01;
		inst_bytes	[490][3]	= 8'h02;
		inst_bytes	[490][4]	= 8'h03;
		inst_bytes	[490][5]	= 8'h04;
		inst_size	[490]		= 4'd6;

		inst_bytes	[491][0]	= 8'h09;
		inst_bytes	[491][1]	= 8'h41;
		inst_bytes	[491][2]	= 8'h01;
		inst_size	[491]		= 4'd3;

		inst_bytes	[492][0]	= 8'h09;
		inst_bytes	[492][1]	= 8'h44;
		inst_bytes	[492][2]	= 8'h52;
		inst_bytes	[492][3]	= 8'h01;
		inst_size	[492]		= 4'd4;

		inst_bytes	[493][0]	= 8'h09;
		inst_bytes	[493][1]	= 8'h81;
		inst_bytes	[493][2]	= 8'h01;
		inst_bytes	[493][3]	= 8'h02;
		inst_bytes	[493][4]	= 8'h03;
		inst_bytes	[493][5]	= 8'h04;
		inst_size	[493]		= 4'd6;

		inst_bytes	[494][0]	= 8'h09;
		inst_bytes	[494][1]	= 8'h84;
		inst_bytes	[494][2]	= 8'h52;
		inst_bytes	[494][3]	= 8'h01;
		inst_bytes	[494][4]	= 8'h02;
		inst_bytes	[494][5]	= 8'h03;
		inst_bytes	[494][6]	= 8'h04;
		inst_size	[494]		= 4'd7;

		inst_bytes	[495][0]	= 8'h09;
		inst_bytes	[495][1]	= 8'hC1;
		inst_size	[495]		= 4'd2;

		inst_bytes	[496][0]	= 8'h0A;
		inst_bytes	[496][1]	= 8'h01;
		inst_size	[496]		= 4'd2;

		inst_bytes	[497][0]	= 8'h0A;
		inst_bytes	[497][1]	= 8'h04;
		inst_bytes	[497][2]	= 8'h52;
		inst_size	[497]		= 4'd3;

		inst_bytes	[498][0]	= 8'h0A;
		inst_bytes	[498][1]	= 8'h05;
		inst_bytes	[498][2]	= 8'h01;
		inst_bytes	[498][3]	= 8'h02;
		inst_bytes	[498][4]	= 8'h03;
		inst_bytes	[498][5]	= 8'h04;
		inst_size	[498]		= 4'd6;

		inst_bytes	[499][0]	= 8'h0A;
		inst_bytes	[499][1]	= 8'h41;
		inst_bytes	[499][2]	= 8'h01;
		inst_size	[499]		= 4'd3;

		inst_bytes	[500][0]	= 8'h0A;
		inst_bytes	[500][1]	= 8'h44;
		inst_bytes	[500][2]	= 8'h52;
		inst_bytes	[500][3]	= 8'h01;
		inst_size	[500]		= 4'd4;

		inst_bytes	[501][0]	= 8'h0A;
		inst_bytes	[501][1]	= 8'h81;
		inst_bytes	[501][2]	= 8'h01;
		inst_bytes	[501][3]	= 8'h02;
		inst_bytes	[501][4]	= 8'h03;
		inst_bytes	[501][5]	= 8'h04;
		inst_size	[501]		= 4'd6;

		inst_bytes	[502][0]	= 8'h0A;
		inst_bytes	[502][1]	= 8'h84;
		inst_bytes	[502][2]	= 8'h52;
		inst_bytes	[502][3]	= 8'h01;
		inst_bytes	[502][4]	= 8'h02;
		inst_bytes	[502][5]	= 8'h03;
		inst_bytes	[502][6]	= 8'h04;
		inst_size	[502]		= 4'd7;

		inst_bytes	[503][0]	= 8'h0A;
		inst_bytes	[503][1]	= 8'hC1;
		inst_size	[503]		= 4'd2;

		inst_bytes	[504][0]	= 8'h0B;
		inst_bytes	[504][1]	= 8'h01;
		inst_size	[504]		= 4'd2;

		inst_bytes	[505][0]	= 8'h0B;
		inst_bytes	[505][1]	= 8'h04;
		inst_bytes	[505][2]	= 8'h52;
		inst_size	[505]		= 4'd3;

		inst_bytes	[506][0]	= 8'h0B;
		inst_bytes	[506][1]	= 8'h05;
		inst_bytes	[506][2]	= 8'h01;
		inst_bytes	[506][3]	= 8'h02;
		inst_bytes	[506][4]	= 8'h03;
		inst_bytes	[506][5]	= 8'h04;
		inst_size	[506]		= 4'd6;

		inst_bytes	[507][0]	= 8'h0B;
		inst_bytes	[507][1]	= 8'h41;
		inst_bytes	[507][2]	= 8'h01;
		inst_size	[507]		= 4'd3;

		inst_bytes	[508][0]	= 8'h0B;
		inst_bytes	[508][1]	= 8'h44;
		inst_bytes	[508][2]	= 8'h52;
		inst_bytes	[508][3]	= 8'h01;
		inst_size	[508]		= 4'd4;

		inst_bytes	[509][0]	= 8'h0B;
		inst_bytes	[509][1]	= 8'h81;
		inst_bytes	[509][2]	= 8'h01;
		inst_bytes	[509][3]	= 8'h02;
		inst_bytes	[509][4]	= 8'h03;
		inst_bytes	[509][5]	= 8'h04;
		inst_size	[509]		= 4'd6;

		inst_bytes	[510][0]	= 8'h0B;
		inst_bytes	[510][1]	= 8'h84;
		inst_bytes	[510][2]	= 8'h52;
		inst_bytes	[510][3]	= 8'h01;
		inst_bytes	[510][4]	= 8'h02;
		inst_bytes	[510][5]	= 8'h03;
		inst_bytes	[510][6]	= 8'h04;
		inst_size	[510]		= 4'd7;

		inst_bytes	[511][0]	= 8'h0B;
		inst_bytes	[511][1]	= 8'hC1;
		inst_size	[511]		= 4'd2;

		inst_bytes	[512][0]	= 8'h0B;
		inst_bytes	[512][1]	= 8'h01;
		inst_size	[512]		= 4'd2;

		inst_bytes	[513][0]	= 8'h0B;
		inst_bytes	[513][1]	= 8'h04;
		inst_bytes	[513][2]	= 8'h52;
		inst_size	[513]		= 4'd3;

		inst_bytes	[514][0]	= 8'h0B;
		inst_bytes	[514][1]	= 8'h05;
		inst_bytes	[514][2]	= 8'h01;
		inst_bytes	[514][3]	= 8'h02;
		inst_bytes	[514][4]	= 8'h03;
		inst_bytes	[514][5]	= 8'h04;
		inst_size	[514]		= 4'd6;

		inst_bytes	[515][0]	= 8'h0B;
		inst_bytes	[515][1]	= 8'h41;
		inst_bytes	[515][2]	= 8'h01;
		inst_size	[515]		= 4'd3;

		inst_bytes	[516][0]	= 8'h0B;
		inst_bytes	[516][1]	= 8'h44;
		inst_bytes	[516][2]	= 8'h52;
		inst_bytes	[516][3]	= 8'h01;
		inst_size	[516]		= 4'd4;

		inst_bytes	[517][0]	= 8'h0B;
		inst_bytes	[517][1]	= 8'h81;
		inst_bytes	[517][2]	= 8'h01;
		inst_bytes	[517][3]	= 8'h02;
		inst_bytes	[517][4]	= 8'h03;
		inst_bytes	[517][5]	= 8'h04;
		inst_size	[517]		= 4'd6;

		inst_bytes	[518][0]	= 8'h0B;
		inst_bytes	[518][1]	= 8'h84;
		inst_bytes	[518][2]	= 8'h52;
		inst_bytes	[518][3]	= 8'h01;
		inst_bytes	[518][4]	= 8'h02;
		inst_bytes	[518][5]	= 8'h03;
		inst_bytes	[518][6]	= 8'h04;
		inst_size	[518]		= 4'd7;

		inst_bytes	[519][0]	= 8'h0B;
		inst_bytes	[519][1]	= 8'hC1;
		inst_size	[519]		= 4'd2;

		inst_bytes	[520][0]	= 8'h0F;
		inst_bytes	[520][1]	= 8'hFD;
		inst_bytes	[520][2]	= 8'h01;
		inst_size	[520]		= 4'd3;

		inst_bytes	[521][0]	= 8'h0F;
		inst_bytes	[521][1]	= 8'hFD;
		inst_bytes	[521][2]	= 8'h04;
		inst_bytes	[521][3]	= 8'h52;
		inst_size	[521]		= 4'd4;

		inst_bytes	[522][0]	= 8'h0F;
		inst_bytes	[522][1]	= 8'hFD;
		inst_bytes	[522][2]	= 8'h05;
		inst_bytes	[522][3]	= 8'h01;
		inst_bytes	[522][4]	= 8'h02;
		inst_bytes	[522][5]	= 8'h03;
		inst_bytes	[522][6]	= 8'h04;
		inst_size	[522]		= 4'd7;

		inst_bytes	[523][0]	= 8'h0F;
		inst_bytes	[523][1]	= 8'hFD;
		inst_bytes	[523][2]	= 8'h41;
		inst_bytes	[523][3]	= 8'h01;
		inst_size	[523]		= 4'd4;

		inst_bytes	[524][0]	= 8'h0F;
		inst_bytes	[524][1]	= 8'hFD;
		inst_bytes	[524][2]	= 8'h44;
		inst_bytes	[524][3]	= 8'h52;
		inst_bytes	[524][4]	= 8'h01;
		inst_size	[524]		= 4'd5;

		inst_bytes	[525][0]	= 8'h0F;
		inst_bytes	[525][1]	= 8'hFD;
		inst_bytes	[525][2]	= 8'h81;
		inst_bytes	[525][3]	= 8'h01;
		inst_bytes	[525][4]	= 8'h02;
		inst_bytes	[525][5]	= 8'h03;
		inst_bytes	[525][6]	= 8'h04;
		inst_size	[525]		= 4'd7;

		inst_bytes	[526][0]	= 8'h0F;
		inst_bytes	[526][1]	= 8'hFD;
		inst_bytes	[526][2]	= 8'h84;
		inst_bytes	[526][3]	= 8'h52;
		inst_bytes	[526][4]	= 8'h01;
		inst_bytes	[526][5]	= 8'h02;
		inst_bytes	[526][6]	= 8'h03;
		inst_bytes	[526][7]	= 8'h04;
		inst_size	[526]		= 4'd8;

		inst_bytes	[527][0]	= 8'h0F;
		inst_bytes	[527][1]	= 8'hFD;
		inst_bytes	[527][2]	= 8'hC1;
		inst_size	[527]		= 4'd3;

		inst_bytes	[528][0]	= 8'h0F;
		inst_bytes	[528][1]	= 8'hFE;
		inst_bytes	[528][2]	= 8'h01;
		inst_size	[528]		= 4'd3;

		inst_bytes	[529][0]	= 8'h0F;
		inst_bytes	[529][1]	= 8'hFE;
		inst_bytes	[529][2]	= 8'h04;
		inst_bytes	[529][3]	= 8'h52;
		inst_size	[529]		= 4'd4;

		inst_bytes	[530][0]	= 8'h0F;
		inst_bytes	[530][1]	= 8'hFE;
		inst_bytes	[530][2]	= 8'h05;
		inst_bytes	[530][3]	= 8'h01;
		inst_bytes	[530][4]	= 8'h02;
		inst_bytes	[530][5]	= 8'h03;
		inst_bytes	[530][6]	= 8'h04;
		inst_size	[530]		= 4'd7;

		inst_bytes	[531][0]	= 8'h0F;
		inst_bytes	[531][1]	= 8'hFE;
		inst_bytes	[531][2]	= 8'h41;
		inst_bytes	[531][3]	= 8'h01;
		inst_size	[531]		= 4'd4;

		inst_bytes	[532][0]	= 8'h0F;
		inst_bytes	[532][1]	= 8'hFE;
		inst_bytes	[532][2]	= 8'h44;
		inst_bytes	[532][3]	= 8'h52;
		inst_bytes	[532][4]	= 8'h01;
		inst_size	[532]		= 4'd5;

		inst_bytes	[533][0]	= 8'h0F;
		inst_bytes	[533][1]	= 8'hFE;
		inst_bytes	[533][2]	= 8'h81;
		inst_bytes	[533][3]	= 8'h01;
		inst_bytes	[533][4]	= 8'h02;
		inst_bytes	[533][5]	= 8'h03;
		inst_bytes	[533][6]	= 8'h04;
		inst_size	[533]		= 4'd7;

		inst_bytes	[534][0]	= 8'h0F;
		inst_bytes	[534][1]	= 8'hFE;
		inst_bytes	[534][2]	= 8'h84;
		inst_bytes	[534][3]	= 8'h52;
		inst_bytes	[534][4]	= 8'h01;
		inst_bytes	[534][5]	= 8'h02;
		inst_bytes	[534][6]	= 8'h03;
		inst_bytes	[534][7]	= 8'h04;
		inst_size	[534]		= 4'd8;

		inst_bytes	[535][0]	= 8'h0F;
		inst_bytes	[535][1]	= 8'hFE;
		inst_bytes	[535][2]	= 8'hC1;
		inst_size	[535]		= 4'd3;

		inst_bytes	[536][0]	= 8'h0F;
		inst_bytes	[536][1]	= 8'hED;
		inst_bytes	[536][2]	= 8'h01;
		inst_size	[536]		= 4'd3;

		inst_bytes	[537][0]	= 8'h0F;
		inst_bytes	[537][1]	= 8'hED;
		inst_bytes	[537][2]	= 8'h04;
		inst_bytes	[537][3]	= 8'h52;
		inst_size	[537]		= 4'd4;

		inst_bytes	[538][0]	= 8'h0F;
		inst_bytes	[538][1]	= 8'hED;
		inst_bytes	[538][2]	= 8'h05;
		inst_bytes	[538][3]	= 8'h01;
		inst_bytes	[538][4]	= 8'h02;
		inst_bytes	[538][5]	= 8'h03;
		inst_bytes	[538][6]	= 8'h04;
		inst_size	[538]		= 4'd7;

		inst_bytes	[539][0]	= 8'h0F;
		inst_bytes	[539][1]	= 8'hED;
		inst_bytes	[539][2]	= 8'h41;
		inst_bytes	[539][3]	= 8'h01;
		inst_size	[539]		= 4'd4;

		inst_bytes	[540][0]	= 8'h0F;
		inst_bytes	[540][1]	= 8'hED;
		inst_bytes	[540][2]	= 8'h44;
		inst_bytes	[540][3]	= 8'h52;
		inst_bytes	[540][4]	= 8'h01;
		inst_size	[540]		= 4'd5;

		inst_bytes	[541][0]	= 8'h0F;
		inst_bytes	[541][1]	= 8'hED;
		inst_bytes	[541][2]	= 8'h81;
		inst_bytes	[541][3]	= 8'h01;
		inst_bytes	[541][4]	= 8'h02;
		inst_bytes	[541][5]	= 8'h03;
		inst_bytes	[541][6]	= 8'h04;
		inst_size	[541]		= 4'd7;

		inst_bytes	[542][0]	= 8'h0F;
		inst_bytes	[542][1]	= 8'hED;
		inst_bytes	[542][2]	= 8'h84;
		inst_bytes	[542][3]	= 8'h52;
		inst_bytes	[542][4]	= 8'h01;
		inst_bytes	[542][5]	= 8'h02;
		inst_bytes	[542][6]	= 8'h03;
		inst_bytes	[542][7]	= 8'h04;
		inst_size	[542]		= 4'd8;

		inst_bytes	[543][0]	= 8'h0F;
		inst_bytes	[543][1]	= 8'hED;
		inst_bytes	[543][2]	= 8'hC1;
		inst_size	[543]		= 4'd3;

		inst_bytes	[544][0]	= 8'h8F;
		inst_bytes	[544][1]	= 8'h01;
		inst_size	[544]		= 4'd2;

		inst_bytes	[545][0]	= 8'h8F;
		inst_bytes	[545][1]	= 8'h04;
		inst_bytes	[545][2]	= 8'h52;
		inst_size	[545]		= 4'd3;

		inst_bytes	[546][0]	= 8'h8F;
		inst_bytes	[546][1]	= 8'h05;
		inst_bytes	[546][2]	= 8'h01;
		inst_bytes	[546][3]	= 8'h02;
		inst_bytes	[546][4]	= 8'h03;
		inst_bytes	[546][5]	= 8'h04;
		inst_size	[546]		= 4'd6;

		inst_bytes	[547][0]	= 8'h8F;
		inst_bytes	[547][1]	= 8'h41;
		inst_bytes	[547][2]	= 8'h01;
		inst_size	[547]		= 4'd3;

		inst_bytes	[548][0]	= 8'h8F;
		inst_bytes	[548][1]	= 8'h44;
		inst_bytes	[548][2]	= 8'h52;
		inst_bytes	[548][3]	= 8'h01;
		inst_size	[548]		= 4'd4;

		inst_bytes	[549][0]	= 8'h8F;
		inst_bytes	[549][1]	= 8'h81;
		inst_bytes	[549][2]	= 8'h01;
		inst_bytes	[549][3]	= 8'h02;
		inst_bytes	[549][4]	= 8'h03;
		inst_bytes	[549][5]	= 8'h04;
		inst_size	[549]		= 4'd6;

		inst_bytes	[550][0]	= 8'h8F;
		inst_bytes	[550][1]	= 8'h84;
		inst_bytes	[550][2]	= 8'h52;
		inst_bytes	[550][3]	= 8'h01;
		inst_bytes	[550][4]	= 8'h02;
		inst_bytes	[550][5]	= 8'h03;
		inst_bytes	[550][6]	= 8'h04;
		inst_size	[550]		= 4'd7;

		inst_bytes	[551][0]	= 8'h8F;
		inst_bytes	[551][1]	= 8'hC1;
		inst_size	[551]		= 4'd2;

		inst_bytes	[552][0]	= 8'h8F;
		inst_bytes	[552][1]	= 8'h01;
		inst_size	[552]		= 4'd2;

		inst_bytes	[553][0]	= 8'h8F;
		inst_bytes	[553][1]	= 8'h04;
		inst_bytes	[553][2]	= 8'h52;
		inst_size	[553]		= 4'd3;

		inst_bytes	[554][0]	= 8'h8F;
		inst_bytes	[554][1]	= 8'h05;
		inst_bytes	[554][2]	= 8'h01;
		inst_bytes	[554][3]	= 8'h02;
		inst_bytes	[554][4]	= 8'h03;
		inst_bytes	[554][5]	= 8'h04;
		inst_size	[554]		= 4'd6;

		inst_bytes	[555][0]	= 8'h8F;
		inst_bytes	[555][1]	= 8'h41;
		inst_bytes	[555][2]	= 8'h01;
		inst_size	[555]		= 4'd3;

		inst_bytes	[556][0]	= 8'h8F;
		inst_bytes	[556][1]	= 8'h44;
		inst_bytes	[556][2]	= 8'h52;
		inst_bytes	[556][3]	= 8'h01;
		inst_size	[556]		= 4'd4;

		inst_bytes	[557][0]	= 8'h8F;
		inst_bytes	[557][1]	= 8'h81;
		inst_bytes	[557][2]	= 8'h01;
		inst_bytes	[557][3]	= 8'h02;
		inst_bytes	[557][4]	= 8'h03;
		inst_bytes	[557][5]	= 8'h04;
		inst_size	[557]		= 4'd6;

		inst_bytes	[558][0]	= 8'h8F;
		inst_bytes	[558][1]	= 8'h84;
		inst_bytes	[558][2]	= 8'h52;
		inst_bytes	[558][3]	= 8'h01;
		inst_bytes	[558][4]	= 8'h02;
		inst_bytes	[558][5]	= 8'h03;
		inst_bytes	[558][6]	= 8'h04;
		inst_size	[558]		= 4'd7;

		inst_bytes	[559][0]	= 8'h8F;
		inst_bytes	[559][1]	= 8'hC1;
		inst_size	[559]		= 4'd2;

		inst_bytes	[560][0]	= 8'h66;
		inst_bytes	[560][1]	= 8'h59;
		inst_size	[560]		= 4'd2;

		inst_bytes	[561][0]	= 8'h59;
		inst_size	[561]		= 4'd1;

		inst_bytes	[562][0]	= 8'h1F;
		inst_size	[562]		= 4'd1;

		inst_bytes	[563][0]	= 8'h07;
		inst_size	[563]		= 4'd1;

		inst_bytes	[564][0]	= 8'h17;
		inst_size	[564]		= 4'd1;

		inst_bytes	[565][0]	= 8'h0F;
		inst_bytes	[565][1]	= 8'hA1;
		inst_size	[565]		= 4'd2;

		inst_bytes	[566][0]	= 8'h0F;
		inst_bytes	[566][1]	= 8'hA9;
		inst_size	[566]		= 4'd2;

		inst_bytes	[567][0]	= 8'h0F;
		inst_bytes	[567][1]	= 8'h70;
		inst_bytes	[567][2]	= 8'h01;
		inst_bytes	[567][3]	= 8'h11;
		inst_size	[567]		= 4'd4;

		inst_bytes	[568][0]	= 8'h0F;
		inst_bytes	[568][1]	= 8'h70;
		inst_bytes	[568][2]	= 8'h04;
		inst_bytes	[568][3]	= 8'h52;
		inst_bytes	[568][4]	= 8'h11;
		inst_size	[568]		= 4'd5;

		inst_bytes	[569][0]	= 8'h0F;
		inst_bytes	[569][1]	= 8'h70;
		inst_bytes	[569][2]	= 8'h05;
		inst_bytes	[569][3]	= 8'h01;
		inst_bytes	[569][4]	= 8'h02;
		inst_bytes	[569][5]	= 8'h03;
		inst_bytes	[569][6]	= 8'h04;
		inst_bytes	[569][7]	= 8'h11;
		inst_size	[569]		= 4'd8;

		inst_bytes	[570][0]	= 8'h0F;
		inst_bytes	[570][1]	= 8'h70;
		inst_bytes	[570][2]	= 8'h41;
		inst_bytes	[570][3]	= 8'h01;
		inst_bytes	[570][4]	= 8'h11;
		inst_size	[570]		= 4'd5;

		inst_bytes	[571][0]	= 8'h0F;
		inst_bytes	[571][1]	= 8'h70;
		inst_bytes	[571][2]	= 8'h44;
		inst_bytes	[571][3]	= 8'h52;
		inst_bytes	[571][4]	= 8'h01;
		inst_bytes	[571][5]	= 8'h11;
		inst_size	[571]		= 4'd6;

		inst_bytes	[572][0]	= 8'h0F;
		inst_bytes	[572][1]	= 8'h70;
		inst_bytes	[572][2]	= 8'h81;
		inst_bytes	[572][3]	= 8'h01;
		inst_bytes	[572][4]	= 8'h02;
		inst_bytes	[572][5]	= 8'h03;
		inst_bytes	[572][6]	= 8'h04;
		inst_bytes	[572][7]	= 8'h11;
		inst_size	[572]		= 4'd8;

		inst_bytes	[573][0]	= 8'h0F;
		inst_bytes	[573][1]	= 8'h70;
		inst_bytes	[573][2]	= 8'h84;
		inst_bytes	[573][3]	= 8'h52;
		inst_bytes	[573][4]	= 8'h01;
		inst_bytes	[573][5]	= 8'h02;
		inst_bytes	[573][6]	= 8'h03;
		inst_bytes	[573][7]	= 8'h04;
		inst_bytes	[573][8]	= 8'h11;
		inst_size	[573]		= 4'd9;

		inst_bytes	[574][0]	= 8'h0F;
		inst_bytes	[574][1]	= 8'h70;
		inst_bytes	[574][2]	= 8'hC1;
		inst_bytes	[574][3]	= 8'h11;
		inst_size	[574]		= 4'd4;

		inst_bytes	[575][0]	= 8'hFF;
		inst_bytes	[575][1]	= 8'h31;
		inst_size	[575]		= 4'd2;

		inst_bytes	[576][0]	= 8'hFF;
		inst_bytes	[576][1]	= 8'h34;
		inst_bytes	[576][2]	= 8'h52;
		inst_size	[576]		= 4'd3;

		inst_bytes	[577][0]	= 8'hFF;
		inst_bytes	[577][1]	= 8'h35;
		inst_bytes	[577][2]	= 8'h01;
		inst_bytes	[577][3]	= 8'h02;
		inst_bytes	[577][4]	= 8'h03;
		inst_bytes	[577][5]	= 8'h04;
		inst_size	[577]		= 4'd6;

		inst_bytes	[578][0]	= 8'hFF;
		inst_bytes	[578][1]	= 8'h71;
		inst_bytes	[578][2]	= 8'h01;
		inst_size	[578]		= 4'd3;

		inst_bytes	[579][0]	= 8'hFF;
		inst_bytes	[579][1]	= 8'h74;
		inst_bytes	[579][2]	= 8'h52;
		inst_bytes	[579][3]	= 8'h01;
		inst_size	[579]		= 4'd4;

		inst_bytes	[580][0]	= 8'hFF;
		inst_bytes	[580][1]	= 8'hB1;
		inst_bytes	[580][2]	= 8'h01;
		inst_bytes	[580][3]	= 8'h02;
		inst_bytes	[580][4]	= 8'h03;
		inst_bytes	[580][5]	= 8'h04;
		inst_size	[580]		= 4'd6;

		inst_bytes	[581][0]	= 8'hFF;
		inst_bytes	[581][1]	= 8'hB4;
		inst_bytes	[581][2]	= 8'h52;
		inst_bytes	[581][3]	= 8'h01;
		inst_bytes	[581][4]	= 8'h02;
		inst_bytes	[581][5]	= 8'h03;
		inst_bytes	[581][6]	= 8'h04;
		inst_size	[581]		= 4'd7;

		inst_bytes	[582][0]	= 8'hFF;
		inst_bytes	[582][1]	= 8'hF1;
		inst_size	[582]		= 4'd2;

		inst_bytes	[583][0]	= 8'hFF;
		inst_bytes	[583][1]	= 8'h31;
		inst_size	[583]		= 4'd2;

		inst_bytes	[584][0]	= 8'hFF;
		inst_bytes	[584][1]	= 8'h34;
		inst_bytes	[584][2]	= 8'h52;
		inst_size	[584]		= 4'd3;

		inst_bytes	[585][0]	= 8'hFF;
		inst_bytes	[585][1]	= 8'h35;
		inst_bytes	[585][2]	= 8'h01;
		inst_bytes	[585][3]	= 8'h02;
		inst_bytes	[585][4]	= 8'h03;
		inst_bytes	[585][5]	= 8'h04;
		inst_size	[585]		= 4'd6;

		inst_bytes	[586][0]	= 8'hFF;
		inst_bytes	[586][1]	= 8'h71;
		inst_bytes	[586][2]	= 8'h01;
		inst_size	[586]		= 4'd3;

		inst_bytes	[587][0]	= 8'hFF;
		inst_bytes	[587][1]	= 8'h74;
		inst_bytes	[587][2]	= 8'h52;
		inst_bytes	[587][3]	= 8'h01;
		inst_size	[587]		= 4'd4;

		inst_bytes	[588][0]	= 8'hFF;
		inst_bytes	[588][1]	= 8'hB1;
		inst_bytes	[588][2]	= 8'h01;
		inst_bytes	[588][3]	= 8'h02;
		inst_bytes	[588][4]	= 8'h03;
		inst_bytes	[588][5]	= 8'h04;
		inst_size	[588]		= 4'd6;

		inst_bytes	[589][0]	= 8'hFF;
		inst_bytes	[589][1]	= 8'hB4;
		inst_bytes	[589][2]	= 8'h52;
		inst_bytes	[589][3]	= 8'h01;
		inst_bytes	[589][4]	= 8'h02;
		inst_bytes	[589][5]	= 8'h03;
		inst_bytes	[589][6]	= 8'h04;
		inst_size	[589]		= 4'd7;

		inst_bytes	[590][0]	= 8'hFF;
		inst_bytes	[590][1]	= 8'hF1;
		inst_size	[590]		= 4'd2;

		inst_bytes	[591][0]	= 8'h66;
		inst_bytes	[591][1]	= 8'h51;
		inst_size	[591]		= 4'd2;

		inst_bytes	[592][0]	= 8'h51;
		inst_size	[592]		= 4'd1;

		inst_bytes	[593][0]	= 8'h6A;
		inst_bytes	[593][1]	= 8'h11;
		inst_size	[593]		= 4'd2;

		inst_bytes	[594][0]	= 8'h66;
		inst_bytes	[594][1]	= 8'h68;
		inst_bytes	[594][2]	= 8'h11;
		inst_bytes	[594][3]	= 8'h12;
		inst_size	[594]		= 4'd4;

		inst_bytes	[595][0]	= 8'h68;
		inst_bytes	[595][1]	= 8'h11;
		inst_bytes	[595][2]	= 8'h12;
		inst_bytes	[595][3]	= 8'h13;
		inst_bytes	[595][4]	= 8'h14;
		inst_size	[595]		= 4'd5;

		inst_bytes	[596][0]	= 8'h0E;
		inst_size	[596]		= 4'd1;

		inst_bytes	[597][0]	= 8'h16;
		inst_size	[597]		= 4'd1;

		inst_bytes	[598][0]	= 8'h1E;
		inst_size	[598]		= 4'd1;

		inst_bytes	[599][0]	= 8'h06;
		inst_size	[599]		= 4'd1;

		inst_bytes	[600][0]	= 8'h0F;
		inst_bytes	[600][1]	= 8'hA0;
		inst_size	[600]		= 4'd2;

		inst_bytes	[601][0]	= 8'h0F;
		inst_bytes	[601][1]	= 8'hA8;
		inst_size	[601]		= 4'd2;

		inst_bytes	[602][0]	= 8'hA6;
		inst_size	[602]		= 4'd1;

		inst_bytes	[603][0]	= 8'hA7;
		inst_size	[603]		= 4'd1;

		inst_bytes	[604][0]	= 8'hA7;
		inst_size	[604]		= 4'd1;

		inst_bytes	[605][0]	= 8'hC3;
		inst_size	[605]		= 4'd1;

		inst_bytes	[606][0]	= 8'hCB;
		inst_size	[606]		= 4'd1;

		inst_bytes	[607][0]	= 8'h66;
		inst_bytes	[607][1]	= 8'hC2;
		inst_bytes	[607][2]	= 8'h11;
		inst_bytes	[607][3]	= 8'h12;
		inst_size	[607]		= 4'd4;

		inst_bytes	[608][0]	= 8'h66;
		inst_bytes	[608][1]	= 8'hCA;
		inst_bytes	[608][2]	= 8'h11;
		inst_bytes	[608][3]	= 8'h12;
		inst_size	[608]		= 4'd4;

		inst_bytes	[609][0]	= 8'hD0;
		inst_bytes	[609][1]	= 8'h21;
		inst_size	[609]		= 4'd2;

		inst_bytes	[610][0]	= 8'hD0;
		inst_bytes	[610][1]	= 8'h24;
		inst_bytes	[610][2]	= 8'h52;
		inst_size	[610]		= 4'd3;

		inst_bytes	[611][0]	= 8'hD0;
		inst_bytes	[611][1]	= 8'h25;
		inst_bytes	[611][2]	= 8'h01;
		inst_bytes	[611][3]	= 8'h02;
		inst_bytes	[611][4]	= 8'h03;
		inst_bytes	[611][5]	= 8'h04;
		inst_size	[611]		= 4'd6;

		inst_bytes	[612][0]	= 8'hD0;
		inst_bytes	[612][1]	= 8'h61;
		inst_bytes	[612][2]	= 8'h01;
		inst_size	[612]		= 4'd3;

		inst_bytes	[613][0]	= 8'hD0;
		inst_bytes	[613][1]	= 8'h64;
		inst_bytes	[613][2]	= 8'h52;
		inst_bytes	[613][3]	= 8'h01;
		inst_size	[613]		= 4'd4;

		inst_bytes	[614][0]	= 8'hD0;
		inst_bytes	[614][1]	= 8'hA1;
		inst_bytes	[614][2]	= 8'h01;
		inst_bytes	[614][3]	= 8'h02;
		inst_bytes	[614][4]	= 8'h03;
		inst_bytes	[614][5]	= 8'h04;
		inst_size	[614]		= 4'd6;

		inst_bytes	[615][0]	= 8'hD0;
		inst_bytes	[615][1]	= 8'hA4;
		inst_bytes	[615][2]	= 8'h52;
		inst_bytes	[615][3]	= 8'h01;
		inst_bytes	[615][4]	= 8'h02;
		inst_bytes	[615][5]	= 8'h03;
		inst_bytes	[615][6]	= 8'h04;
		inst_size	[615]		= 4'd7;

		inst_bytes	[616][0]	= 8'hD0;
		inst_bytes	[616][1]	= 8'hE1;
		inst_size	[616]		= 4'd2;

		inst_bytes	[617][0]	= 8'hD2;
		inst_bytes	[617][1]	= 8'h21;
		inst_size	[617]		= 4'd2;

		inst_bytes	[618][0]	= 8'hD2;
		inst_bytes	[618][1]	= 8'h24;
		inst_bytes	[618][2]	= 8'h52;
		inst_size	[618]		= 4'd3;

		inst_bytes	[619][0]	= 8'hD2;
		inst_bytes	[619][1]	= 8'h25;
		inst_bytes	[619][2]	= 8'h01;
		inst_bytes	[619][3]	= 8'h02;
		inst_bytes	[619][4]	= 8'h03;
		inst_bytes	[619][5]	= 8'h04;
		inst_size	[619]		= 4'd6;

		inst_bytes	[620][0]	= 8'hD2;
		inst_bytes	[620][1]	= 8'h61;
		inst_bytes	[620][2]	= 8'h01;
		inst_size	[620]		= 4'd3;

		inst_bytes	[621][0]	= 8'hD2;
		inst_bytes	[621][1]	= 8'h64;
		inst_bytes	[621][2]	= 8'h52;
		inst_bytes	[621][3]	= 8'h01;
		inst_size	[621]		= 4'd4;

		inst_bytes	[622][0]	= 8'hD2;
		inst_bytes	[622][1]	= 8'hA1;
		inst_bytes	[622][2]	= 8'h01;
		inst_bytes	[622][3]	= 8'h02;
		inst_bytes	[622][4]	= 8'h03;
		inst_bytes	[622][5]	= 8'h04;
		inst_size	[622]		= 4'd6;

		inst_bytes	[623][0]	= 8'hD2;
		inst_bytes	[623][1]	= 8'hA4;
		inst_bytes	[623][2]	= 8'h52;
		inst_bytes	[623][3]	= 8'h01;
		inst_bytes	[623][4]	= 8'h02;
		inst_bytes	[623][5]	= 8'h03;
		inst_bytes	[623][6]	= 8'h04;
		inst_size	[623]		= 4'd7;

		inst_bytes	[624][0]	= 8'hD2;
		inst_bytes	[624][1]	= 8'hE1;
		inst_size	[624]		= 4'd2;

		inst_bytes	[625][0]	= 8'hC0;
		inst_bytes	[625][1]	= 8'h21;
		inst_bytes	[625][2]	= 8'h11;
		inst_size	[625]		= 4'd3;

		inst_bytes	[626][0]	= 8'hC0;
		inst_bytes	[626][1]	= 8'h24;
		inst_bytes	[626][2]	= 8'h52;
		inst_bytes	[626][3]	= 8'h11;
		inst_size	[626]		= 4'd4;

		inst_bytes	[627][0]	= 8'hC0;
		inst_bytes	[627][1]	= 8'h25;
		inst_bytes	[627][2]	= 8'h01;
		inst_bytes	[627][3]	= 8'h02;
		inst_bytes	[627][4]	= 8'h03;
		inst_bytes	[627][5]	= 8'h04;
		inst_bytes	[627][6]	= 8'h11;
		inst_size	[627]		= 4'd7;

		inst_bytes	[628][0]	= 8'hC0;
		inst_bytes	[628][1]	= 8'h61;
		inst_bytes	[628][2]	= 8'h01;
		inst_bytes	[628][3]	= 8'h11;
		inst_size	[628]		= 4'd4;

		inst_bytes	[629][0]	= 8'hC0;
		inst_bytes	[629][1]	= 8'h64;
		inst_bytes	[629][2]	= 8'h52;
		inst_bytes	[629][3]	= 8'h01;
		inst_bytes	[629][4]	= 8'h11;
		inst_size	[629]		= 4'd5;

		inst_bytes	[630][0]	= 8'hC0;
		inst_bytes	[630][1]	= 8'hA1;
		inst_bytes	[630][2]	= 8'h01;
		inst_bytes	[630][3]	= 8'h02;
		inst_bytes	[630][4]	= 8'h03;
		inst_bytes	[630][5]	= 8'h04;
		inst_bytes	[630][6]	= 8'h11;
		inst_size	[630]		= 4'd7;

		inst_bytes	[631][0]	= 8'hC0;
		inst_bytes	[631][1]	= 8'hA4;
		inst_bytes	[631][2]	= 8'h52;
		inst_bytes	[631][3]	= 8'h01;
		inst_bytes	[631][4]	= 8'h02;
		inst_bytes	[631][5]	= 8'h03;
		inst_bytes	[631][6]	= 8'h04;
		inst_bytes	[631][7]	= 8'h11;
		inst_size	[631]		= 4'd8;

		inst_bytes	[632][0]	= 8'hC0;
		inst_bytes	[632][1]	= 8'hE1;
		inst_bytes	[632][2]	= 8'h11;
		inst_size	[632]		= 4'd3;

		inst_bytes	[633][0]	= 8'hD1;
		inst_bytes	[633][1]	= 8'h21;
		inst_size	[633]		= 4'd2;

		inst_bytes	[634][0]	= 8'hD1;
		inst_bytes	[634][1]	= 8'h24;
		inst_bytes	[634][2]	= 8'h52;
		inst_size	[634]		= 4'd3;

		inst_bytes	[635][0]	= 8'hD1;
		inst_bytes	[635][1]	= 8'h25;
		inst_bytes	[635][2]	= 8'h01;
		inst_bytes	[635][3]	= 8'h02;
		inst_bytes	[635][4]	= 8'h03;
		inst_bytes	[635][5]	= 8'h04;
		inst_size	[635]		= 4'd6;

		inst_bytes	[636][0]	= 8'hD1;
		inst_bytes	[636][1]	= 8'h61;
		inst_bytes	[636][2]	= 8'h01;
		inst_size	[636]		= 4'd3;

		inst_bytes	[637][0]	= 8'hD1;
		inst_bytes	[637][1]	= 8'h64;
		inst_bytes	[637][2]	= 8'h52;
		inst_bytes	[637][3]	= 8'h01;
		inst_size	[637]		= 4'd4;

		inst_bytes	[638][0]	= 8'hD1;
		inst_bytes	[638][1]	= 8'hA1;
		inst_bytes	[638][2]	= 8'h01;
		inst_bytes	[638][3]	= 8'h02;
		inst_bytes	[638][4]	= 8'h03;
		inst_bytes	[638][5]	= 8'h04;
		inst_size	[638]		= 4'd6;

		inst_bytes	[639][0]	= 8'hD1;
		inst_bytes	[639][1]	= 8'hA4;
		inst_bytes	[639][2]	= 8'h52;
		inst_bytes	[639][3]	= 8'h01;
		inst_bytes	[639][4]	= 8'h02;
		inst_bytes	[639][5]	= 8'h03;
		inst_bytes	[639][6]	= 8'h04;
		inst_size	[639]		= 4'd7;

		inst_bytes	[640][0]	= 8'hD1;
		inst_bytes	[640][1]	= 8'hE1;
		inst_size	[640]		= 4'd2;

		inst_bytes	[641][0]	= 8'hD3;
		inst_bytes	[641][1]	= 8'h21;
		inst_size	[641]		= 4'd2;

		inst_bytes	[642][0]	= 8'hD3;
		inst_bytes	[642][1]	= 8'h24;
		inst_bytes	[642][2]	= 8'h52;
		inst_size	[642]		= 4'd3;

		inst_bytes	[643][0]	= 8'hD3;
		inst_bytes	[643][1]	= 8'h25;
		inst_bytes	[643][2]	= 8'h01;
		inst_bytes	[643][3]	= 8'h02;
		inst_bytes	[643][4]	= 8'h03;
		inst_bytes	[643][5]	= 8'h04;
		inst_size	[643]		= 4'd6;

		inst_bytes	[644][0]	= 8'hD3;
		inst_bytes	[644][1]	= 8'h61;
		inst_bytes	[644][2]	= 8'h01;
		inst_size	[644]		= 4'd3;

		inst_bytes	[645][0]	= 8'hD3;
		inst_bytes	[645][1]	= 8'h64;
		inst_bytes	[645][2]	= 8'h52;
		inst_bytes	[645][3]	= 8'h01;
		inst_size	[645]		= 4'd4;

		inst_bytes	[646][0]	= 8'hD3;
		inst_bytes	[646][1]	= 8'hA1;
		inst_bytes	[646][2]	= 8'h01;
		inst_bytes	[646][3]	= 8'h02;
		inst_bytes	[646][4]	= 8'h03;
		inst_bytes	[646][5]	= 8'h04;
		inst_size	[646]		= 4'd6;

		inst_bytes	[647][0]	= 8'hD3;
		inst_bytes	[647][1]	= 8'hA4;
		inst_bytes	[647][2]	= 8'h52;
		inst_bytes	[647][3]	= 8'h01;
		inst_bytes	[647][4]	= 8'h02;
		inst_bytes	[647][5]	= 8'h03;
		inst_bytes	[647][6]	= 8'h04;
		inst_size	[647]		= 4'd7;

		inst_bytes	[648][0]	= 8'hD3;
		inst_bytes	[648][1]	= 8'hE1;
		inst_size	[648]		= 4'd2;

		inst_bytes	[649][0]	= 8'hC1;
		inst_bytes	[649][1]	= 8'h21;
		inst_bytes	[649][2]	= 8'h11;
		inst_size	[649]		= 4'd3;

		inst_bytes	[650][0]	= 8'hC1;
		inst_bytes	[650][1]	= 8'h24;
		inst_bytes	[650][2]	= 8'h52;
		inst_bytes	[650][3]	= 8'h11;
		inst_size	[650]		= 4'd4;

		inst_bytes	[651][0]	= 8'hC1;
		inst_bytes	[651][1]	= 8'h25;
		inst_bytes	[651][2]	= 8'h01;
		inst_bytes	[651][3]	= 8'h02;
		inst_bytes	[651][4]	= 8'h03;
		inst_bytes	[651][5]	= 8'h04;
		inst_bytes	[651][6]	= 8'h11;
		inst_size	[651]		= 4'd7;

		inst_bytes	[652][0]	= 8'hC1;
		inst_bytes	[652][1]	= 8'h61;
		inst_bytes	[652][2]	= 8'h01;
		inst_bytes	[652][3]	= 8'h11;
		inst_size	[652]		= 4'd4;

		inst_bytes	[653][0]	= 8'hC1;
		inst_bytes	[653][1]	= 8'h64;
		inst_bytes	[653][2]	= 8'h52;
		inst_bytes	[653][3]	= 8'h01;
		inst_bytes	[653][4]	= 8'h11;
		inst_size	[653]		= 4'd5;

		inst_bytes	[654][0]	= 8'hC1;
		inst_bytes	[654][1]	= 8'hA1;
		inst_bytes	[654][2]	= 8'h01;
		inst_bytes	[654][3]	= 8'h02;
		inst_bytes	[654][4]	= 8'h03;
		inst_bytes	[654][5]	= 8'h04;
		inst_bytes	[654][6]	= 8'h11;
		inst_size	[654]		= 4'd7;

		inst_bytes	[655][0]	= 8'hC1;
		inst_bytes	[655][1]	= 8'hA4;
		inst_bytes	[655][2]	= 8'h52;
		inst_bytes	[655][3]	= 8'h01;
		inst_bytes	[655][4]	= 8'h02;
		inst_bytes	[655][5]	= 8'h03;
		inst_bytes	[655][6]	= 8'h04;
		inst_bytes	[655][7]	= 8'h11;
		inst_size	[655]		= 4'd8;

		inst_bytes	[656][0]	= 8'hC1;
		inst_bytes	[656][1]	= 8'hE1;
		inst_bytes	[656][2]	= 8'h11;
		inst_size	[656]		= 4'd3;

		inst_bytes	[657][0]	= 8'hD1;
		inst_bytes	[657][1]	= 8'h21;
		inst_size	[657]		= 4'd2;

		inst_bytes	[658][0]	= 8'hD1;
		inst_bytes	[658][1]	= 8'h24;
		inst_bytes	[658][2]	= 8'h52;
		inst_size	[658]		= 4'd3;

		inst_bytes	[659][0]	= 8'hD1;
		inst_bytes	[659][1]	= 8'h25;
		inst_bytes	[659][2]	= 8'h01;
		inst_bytes	[659][3]	= 8'h02;
		inst_bytes	[659][4]	= 8'h03;
		inst_bytes	[659][5]	= 8'h04;
		inst_size	[659]		= 4'd6;

		inst_bytes	[660][0]	= 8'hD1;
		inst_bytes	[660][1]	= 8'h61;
		inst_bytes	[660][2]	= 8'h01;
		inst_size	[660]		= 4'd3;

		inst_bytes	[661][0]	= 8'hD1;
		inst_bytes	[661][1]	= 8'h64;
		inst_bytes	[661][2]	= 8'h52;
		inst_bytes	[661][3]	= 8'h01;
		inst_size	[661]		= 4'd4;

		inst_bytes	[662][0]	= 8'hD1;
		inst_bytes	[662][1]	= 8'hA1;
		inst_bytes	[662][2]	= 8'h01;
		inst_bytes	[662][3]	= 8'h02;
		inst_bytes	[662][4]	= 8'h03;
		inst_bytes	[662][5]	= 8'h04;
		inst_size	[662]		= 4'd6;

		inst_bytes	[663][0]	= 8'hD1;
		inst_bytes	[663][1]	= 8'hA4;
		inst_bytes	[663][2]	= 8'h52;
		inst_bytes	[663][3]	= 8'h01;
		inst_bytes	[663][4]	= 8'h02;
		inst_bytes	[663][5]	= 8'h03;
		inst_bytes	[663][6]	= 8'h04;
		inst_size	[663]		= 4'd7;

		inst_bytes	[664][0]	= 8'hD1;
		inst_bytes	[664][1]	= 8'hE1;
		inst_size	[664]		= 4'd2;

		inst_bytes	[665][0]	= 8'hD3;
		inst_bytes	[665][1]	= 8'h21;
		inst_size	[665]		= 4'd2;

		inst_bytes	[666][0]	= 8'hD3;
		inst_bytes	[666][1]	= 8'h24;
		inst_bytes	[666][2]	= 8'h52;
		inst_size	[666]		= 4'd3;

		inst_bytes	[667][0]	= 8'hD3;
		inst_bytes	[667][1]	= 8'h25;
		inst_bytes	[667][2]	= 8'h01;
		inst_bytes	[667][3]	= 8'h02;
		inst_bytes	[667][4]	= 8'h03;
		inst_bytes	[667][5]	= 8'h04;
		inst_size	[667]		= 4'd6;

		inst_bytes	[668][0]	= 8'hD3;
		inst_bytes	[668][1]	= 8'h61;
		inst_bytes	[668][2]	= 8'h01;
		inst_size	[668]		= 4'd3;

		inst_bytes	[669][0]	= 8'hD3;
		inst_bytes	[669][1]	= 8'h64;
		inst_bytes	[669][2]	= 8'h52;
		inst_bytes	[669][3]	= 8'h01;
		inst_size	[669]		= 4'd4;

		inst_bytes	[670][0]	= 8'hD3;
		inst_bytes	[670][1]	= 8'hA1;
		inst_bytes	[670][2]	= 8'h01;
		inst_bytes	[670][3]	= 8'h02;
		inst_bytes	[670][4]	= 8'h03;
		inst_bytes	[670][5]	= 8'h04;
		inst_size	[670]		= 4'd6;

		inst_bytes	[671][0]	= 8'hD3;
		inst_bytes	[671][1]	= 8'hA4;
		inst_bytes	[671][2]	= 8'h52;
		inst_bytes	[671][3]	= 8'h01;
		inst_bytes	[671][4]	= 8'h02;
		inst_bytes	[671][5]	= 8'h03;
		inst_bytes	[671][6]	= 8'h04;
		inst_size	[671]		= 4'd7;

		inst_bytes	[672][0]	= 8'hD3;
		inst_bytes	[672][1]	= 8'hE1;
		inst_size	[672]		= 4'd2;

		inst_bytes	[673][0]	= 8'hC1;
		inst_bytes	[673][1]	= 8'h21;
		inst_bytes	[673][2]	= 8'h11;
		inst_size	[673]		= 4'd3;

		inst_bytes	[674][0]	= 8'hC1;
		inst_bytes	[674][1]	= 8'h24;
		inst_bytes	[674][2]	= 8'h52;
		inst_bytes	[674][3]	= 8'h11;
		inst_size	[674]		= 4'd4;

		inst_bytes	[675][0]	= 8'hC1;
		inst_bytes	[675][1]	= 8'h25;
		inst_bytes	[675][2]	= 8'h01;
		inst_bytes	[675][3]	= 8'h02;
		inst_bytes	[675][4]	= 8'h03;
		inst_bytes	[675][5]	= 8'h04;
		inst_bytes	[675][6]	= 8'h11;
		inst_size	[675]		= 4'd7;

		inst_bytes	[676][0]	= 8'hC1;
		inst_bytes	[676][1]	= 8'h61;
		inst_bytes	[676][2]	= 8'h01;
		inst_bytes	[676][3]	= 8'h11;
		inst_size	[676]		= 4'd4;

		inst_bytes	[677][0]	= 8'hC1;
		inst_bytes	[677][1]	= 8'h64;
		inst_bytes	[677][2]	= 8'h52;
		inst_bytes	[677][3]	= 8'h01;
		inst_bytes	[677][4]	= 8'h11;
		inst_size	[677]		= 4'd5;

		inst_bytes	[678][0]	= 8'hC1;
		inst_bytes	[678][1]	= 8'hA1;
		inst_bytes	[678][2]	= 8'h01;
		inst_bytes	[678][3]	= 8'h02;
		inst_bytes	[678][4]	= 8'h03;
		inst_bytes	[678][5]	= 8'h04;
		inst_bytes	[678][6]	= 8'h11;
		inst_size	[678]		= 4'd7;

		inst_bytes	[679][0]	= 8'hC1;
		inst_bytes	[679][1]	= 8'hA4;
		inst_bytes	[679][2]	= 8'h52;
		inst_bytes	[679][3]	= 8'h01;
		inst_bytes	[679][4]	= 8'h02;
		inst_bytes	[679][5]	= 8'h03;
		inst_bytes	[679][6]	= 8'h04;
		inst_bytes	[679][7]	= 8'h11;
		inst_size	[679]		= 4'd8;

		inst_bytes	[680][0]	= 8'hC1;
		inst_bytes	[680][1]	= 8'hE1;
		inst_bytes	[680][2]	= 8'h11;
		inst_size	[680]		= 4'd3;

		inst_bytes	[681][0]	= 8'hD0;
		inst_bytes	[681][1]	= 8'h39;
		inst_size	[681]		= 4'd2;

		inst_bytes	[682][0]	= 8'hD0;
		inst_bytes	[682][1]	= 8'h3C;
		inst_bytes	[682][2]	= 8'h52;
		inst_size	[682]		= 4'd3;

		inst_bytes	[683][0]	= 8'hD0;
		inst_bytes	[683][1]	= 8'h3D;
		inst_bytes	[683][2]	= 8'h01;
		inst_bytes	[683][3]	= 8'h02;
		inst_bytes	[683][4]	= 8'h03;
		inst_bytes	[683][5]	= 8'h04;
		inst_size	[683]		= 4'd6;

		inst_bytes	[684][0]	= 8'hD0;
		inst_bytes	[684][1]	= 8'h79;
		inst_bytes	[684][2]	= 8'h01;
		inst_size	[684]		= 4'd3;

		inst_bytes	[685][0]	= 8'hD0;
		inst_bytes	[685][1]	= 8'h7C;
		inst_bytes	[685][2]	= 8'h52;
		inst_bytes	[685][3]	= 8'h01;
		inst_size	[685]		= 4'd4;

		inst_bytes	[686][0]	= 8'hD0;
		inst_bytes	[686][1]	= 8'hB9;
		inst_bytes	[686][2]	= 8'h01;
		inst_bytes	[686][3]	= 8'h02;
		inst_bytes	[686][4]	= 8'h03;
		inst_bytes	[686][5]	= 8'h04;
		inst_size	[686]		= 4'd6;

		inst_bytes	[687][0]	= 8'hD0;
		inst_bytes	[687][1]	= 8'hBC;
		inst_bytes	[687][2]	= 8'h52;
		inst_bytes	[687][3]	= 8'h01;
		inst_bytes	[687][4]	= 8'h02;
		inst_bytes	[687][5]	= 8'h03;
		inst_bytes	[687][6]	= 8'h04;
		inst_size	[687]		= 4'd7;

		inst_bytes	[688][0]	= 8'hD0;
		inst_bytes	[688][1]	= 8'hF9;
		inst_size	[688]		= 4'd2;

		inst_bytes	[689][0]	= 8'hD2;
		inst_bytes	[689][1]	= 8'h39;
		inst_size	[689]		= 4'd2;

		inst_bytes	[690][0]	= 8'hD2;
		inst_bytes	[690][1]	= 8'h3C;
		inst_bytes	[690][2]	= 8'h52;
		inst_size	[690]		= 4'd3;

		inst_bytes	[691][0]	= 8'hD2;
		inst_bytes	[691][1]	= 8'h3D;
		inst_bytes	[691][2]	= 8'h01;
		inst_bytes	[691][3]	= 8'h02;
		inst_bytes	[691][4]	= 8'h03;
		inst_bytes	[691][5]	= 8'h04;
		inst_size	[691]		= 4'd6;

		inst_bytes	[692][0]	= 8'hD2;
		inst_bytes	[692][1]	= 8'h79;
		inst_bytes	[692][2]	= 8'h01;
		inst_size	[692]		= 4'd3;

		inst_bytes	[693][0]	= 8'hD2;
		inst_bytes	[693][1]	= 8'h7C;
		inst_bytes	[693][2]	= 8'h52;
		inst_bytes	[693][3]	= 8'h01;
		inst_size	[693]		= 4'd4;

		inst_bytes	[694][0]	= 8'hD2;
		inst_bytes	[694][1]	= 8'hB9;
		inst_bytes	[694][2]	= 8'h01;
		inst_bytes	[694][3]	= 8'h02;
		inst_bytes	[694][4]	= 8'h03;
		inst_bytes	[694][5]	= 8'h04;
		inst_size	[694]		= 4'd6;

		inst_bytes	[695][0]	= 8'hD2;
		inst_bytes	[695][1]	= 8'hBC;
		inst_bytes	[695][2]	= 8'h52;
		inst_bytes	[695][3]	= 8'h01;
		inst_bytes	[695][4]	= 8'h02;
		inst_bytes	[695][5]	= 8'h03;
		inst_bytes	[695][6]	= 8'h04;
		inst_size	[695]		= 4'd7;

		inst_bytes	[696][0]	= 8'hD2;
		inst_bytes	[696][1]	= 8'hF9;
		inst_size	[696]		= 4'd2;

		inst_bytes	[697][0]	= 8'hC0;
		inst_bytes	[697][1]	= 8'h39;
		inst_bytes	[697][2]	= 8'h11;
		inst_size	[697]		= 4'd3;

		inst_bytes	[698][0]	= 8'hC0;
		inst_bytes	[698][1]	= 8'h3C;
		inst_bytes	[698][2]	= 8'h52;
		inst_bytes	[698][3]	= 8'h11;
		inst_size	[698]		= 4'd4;

		inst_bytes	[699][0]	= 8'hC0;
		inst_bytes	[699][1]	= 8'h3D;
		inst_bytes	[699][2]	= 8'h01;
		inst_bytes	[699][3]	= 8'h02;
		inst_bytes	[699][4]	= 8'h03;
		inst_bytes	[699][5]	= 8'h04;
		inst_bytes	[699][6]	= 8'h11;
		inst_size	[699]		= 4'd7;

		inst_bytes	[700][0]	= 8'hC0;
		inst_bytes	[700][1]	= 8'h79;
		inst_bytes	[700][2]	= 8'h01;
		inst_bytes	[700][3]	= 8'h11;
		inst_size	[700]		= 4'd4;

		inst_bytes	[701][0]	= 8'hC0;
		inst_bytes	[701][1]	= 8'h7C;
		inst_bytes	[701][2]	= 8'h52;
		inst_bytes	[701][3]	= 8'h01;
		inst_bytes	[701][4]	= 8'h11;
		inst_size	[701]		= 4'd5;

		inst_bytes	[702][0]	= 8'hC0;
		inst_bytes	[702][1]	= 8'hB9;
		inst_bytes	[702][2]	= 8'h01;
		inst_bytes	[702][3]	= 8'h02;
		inst_bytes	[702][4]	= 8'h03;
		inst_bytes	[702][5]	= 8'h04;
		inst_bytes	[702][6]	= 8'h11;
		inst_size	[702]		= 4'd7;

		inst_bytes	[703][0]	= 8'hC0;
		inst_bytes	[703][1]	= 8'hBC;
		inst_bytes	[703][2]	= 8'h52;
		inst_bytes	[703][3]	= 8'h01;
		inst_bytes	[703][4]	= 8'h02;
		inst_bytes	[703][5]	= 8'h03;
		inst_bytes	[703][6]	= 8'h04;
		inst_bytes	[703][7]	= 8'h11;
		inst_size	[703]		= 4'd8;

		inst_bytes	[704][0]	= 8'hC0;
		inst_bytes	[704][1]	= 8'hF9;
		inst_bytes	[704][2]	= 8'h11;
		inst_size	[704]		= 4'd3;

		inst_bytes	[705][0]	= 8'hD1;
		inst_bytes	[705][1]	= 8'h39;
		inst_size	[705]		= 4'd2;

		inst_bytes	[706][0]	= 8'hD1;
		inst_bytes	[706][1]	= 8'h3C;
		inst_bytes	[706][2]	= 8'h52;
		inst_size	[706]		= 4'd3;

		inst_bytes	[707][0]	= 8'hD1;
		inst_bytes	[707][1]	= 8'h3D;
		inst_bytes	[707][2]	= 8'h01;
		inst_bytes	[707][3]	= 8'h02;
		inst_bytes	[707][4]	= 8'h03;
		inst_bytes	[707][5]	= 8'h04;
		inst_size	[707]		= 4'd6;

		inst_bytes	[708][0]	= 8'hD1;
		inst_bytes	[708][1]	= 8'h79;
		inst_bytes	[708][2]	= 8'h01;
		inst_size	[708]		= 4'd3;

		inst_bytes	[709][0]	= 8'hD1;
		inst_bytes	[709][1]	= 8'h7C;
		inst_bytes	[709][2]	= 8'h52;
		inst_bytes	[709][3]	= 8'h01;
		inst_size	[709]		= 4'd4;

		inst_bytes	[710][0]	= 8'hD1;
		inst_bytes	[710][1]	= 8'hB9;
		inst_bytes	[710][2]	= 8'h01;
		inst_bytes	[710][3]	= 8'h02;
		inst_bytes	[710][4]	= 8'h03;
		inst_bytes	[710][5]	= 8'h04;
		inst_size	[710]		= 4'd6;

		inst_bytes	[711][0]	= 8'hD1;
		inst_bytes	[711][1]	= 8'hBC;
		inst_bytes	[711][2]	= 8'h52;
		inst_bytes	[711][3]	= 8'h01;
		inst_bytes	[711][4]	= 8'h02;
		inst_bytes	[711][5]	= 8'h03;
		inst_bytes	[711][6]	= 8'h04;
		inst_size	[711]		= 4'd7;

		inst_bytes	[712][0]	= 8'hD1;
		inst_bytes	[712][1]	= 8'hF9;
		inst_size	[712]		= 4'd2;

		inst_bytes	[713][0]	= 8'hD3;
		inst_bytes	[713][1]	= 8'h39;
		inst_size	[713]		= 4'd2;

		inst_bytes	[714][0]	= 8'hD3;
		inst_bytes	[714][1]	= 8'h3C;
		inst_bytes	[714][2]	= 8'h52;
		inst_size	[714]		= 4'd3;

		inst_bytes	[715][0]	= 8'hD3;
		inst_bytes	[715][1]	= 8'h3D;
		inst_bytes	[715][2]	= 8'h01;
		inst_bytes	[715][3]	= 8'h02;
		inst_bytes	[715][4]	= 8'h03;
		inst_bytes	[715][5]	= 8'h04;
		inst_size	[715]		= 4'd6;

		inst_bytes	[716][0]	= 8'hD3;
		inst_bytes	[716][1]	= 8'h79;
		inst_bytes	[716][2]	= 8'h01;
		inst_size	[716]		= 4'd3;

		inst_bytes	[717][0]	= 8'hD3;
		inst_bytes	[717][1]	= 8'h7C;
		inst_bytes	[717][2]	= 8'h52;
		inst_bytes	[717][3]	= 8'h01;
		inst_size	[717]		= 4'd4;

		inst_bytes	[718][0]	= 8'hD3;
		inst_bytes	[718][1]	= 8'hB9;
		inst_bytes	[718][2]	= 8'h01;
		inst_bytes	[718][3]	= 8'h02;
		inst_bytes	[718][4]	= 8'h03;
		inst_bytes	[718][5]	= 8'h04;
		inst_size	[718]		= 4'd6;

		inst_bytes	[719][0]	= 8'hD3;
		inst_bytes	[719][1]	= 8'hBC;
		inst_bytes	[719][2]	= 8'h52;
		inst_bytes	[719][3]	= 8'h01;
		inst_bytes	[719][4]	= 8'h02;
		inst_bytes	[719][5]	= 8'h03;
		inst_bytes	[719][6]	= 8'h04;
		inst_size	[719]		= 4'd7;

		inst_bytes	[720][0]	= 8'hD3;
		inst_bytes	[720][1]	= 8'hF9;
		inst_size	[720]		= 4'd2;

		inst_bytes	[721][0]	= 8'hC1;
		inst_bytes	[721][1]	= 8'h39;
		inst_bytes	[721][2]	= 8'h11;
		inst_size	[721]		= 4'd3;

		inst_bytes	[722][0]	= 8'hC1;
		inst_bytes	[722][1]	= 8'h3C;
		inst_bytes	[722][2]	= 8'h52;
		inst_bytes	[722][3]	= 8'h11;
		inst_size	[722]		= 4'd4;

		inst_bytes	[723][0]	= 8'hC1;
		inst_bytes	[723][1]	= 8'h3D;
		inst_bytes	[723][2]	= 8'h01;
		inst_bytes	[723][3]	= 8'h02;
		inst_bytes	[723][4]	= 8'h03;
		inst_bytes	[723][5]	= 8'h04;
		inst_bytes	[723][6]	= 8'h11;
		inst_size	[723]		= 4'd7;

		inst_bytes	[724][0]	= 8'hC1;
		inst_bytes	[724][1]	= 8'h79;
		inst_bytes	[724][2]	= 8'h01;
		inst_bytes	[724][3]	= 8'h11;
		inst_size	[724]		= 4'd4;

		inst_bytes	[725][0]	= 8'hC1;
		inst_bytes	[725][1]	= 8'h7C;
		inst_bytes	[725][2]	= 8'h52;
		inst_bytes	[725][3]	= 8'h01;
		inst_bytes	[725][4]	= 8'h11;
		inst_size	[725]		= 4'd5;

		inst_bytes	[726][0]	= 8'hC1;
		inst_bytes	[726][1]	= 8'hB9;
		inst_bytes	[726][2]	= 8'h01;
		inst_bytes	[726][3]	= 8'h02;
		inst_bytes	[726][4]	= 8'h03;
		inst_bytes	[726][5]	= 8'h04;
		inst_bytes	[726][6]	= 8'h11;
		inst_size	[726]		= 4'd7;

		inst_bytes	[727][0]	= 8'hC1;
		inst_bytes	[727][1]	= 8'hBC;
		inst_bytes	[727][2]	= 8'h52;
		inst_bytes	[727][3]	= 8'h01;
		inst_bytes	[727][4]	= 8'h02;
		inst_bytes	[727][5]	= 8'h03;
		inst_bytes	[727][6]	= 8'h04;
		inst_bytes	[727][7]	= 8'h11;
		inst_size	[727]		= 4'd8;

		inst_bytes	[728][0]	= 8'hC1;
		inst_bytes	[728][1]	= 8'hF9;
		inst_bytes	[728][2]	= 8'h11;
		inst_size	[728]		= 4'd3;

		inst_bytes	[729][0]	= 8'hD1;
		inst_bytes	[729][1]	= 8'h39;
		inst_size	[729]		= 4'd2;

		inst_bytes	[730][0]	= 8'hD1;
		inst_bytes	[730][1]	= 8'h3C;
		inst_bytes	[730][2]	= 8'h52;
		inst_size	[730]		= 4'd3;

		inst_bytes	[731][0]	= 8'hD1;
		inst_bytes	[731][1]	= 8'h3D;
		inst_bytes	[731][2]	= 8'h01;
		inst_bytes	[731][3]	= 8'h02;
		inst_bytes	[731][4]	= 8'h03;
		inst_bytes	[731][5]	= 8'h04;
		inst_size	[731]		= 4'd6;

		inst_bytes	[732][0]	= 8'hD1;
		inst_bytes	[732][1]	= 8'h79;
		inst_bytes	[732][2]	= 8'h01;
		inst_size	[732]		= 4'd3;

		inst_bytes	[733][0]	= 8'hD1;
		inst_bytes	[733][1]	= 8'h7C;
		inst_bytes	[733][2]	= 8'h52;
		inst_bytes	[733][3]	= 8'h01;
		inst_size	[733]		= 4'd4;

		inst_bytes	[734][0]	= 8'hD1;
		inst_bytes	[734][1]	= 8'hB9;
		inst_bytes	[734][2]	= 8'h01;
		inst_bytes	[734][3]	= 8'h02;
		inst_bytes	[734][4]	= 8'h03;
		inst_bytes	[734][5]	= 8'h04;
		inst_size	[734]		= 4'd6;

		inst_bytes	[735][0]	= 8'hD1;
		inst_bytes	[735][1]	= 8'hBC;
		inst_bytes	[735][2]	= 8'h52;
		inst_bytes	[735][3]	= 8'h01;
		inst_bytes	[735][4]	= 8'h02;
		inst_bytes	[735][5]	= 8'h03;
		inst_bytes	[735][6]	= 8'h04;
		inst_size	[735]		= 4'd7;

		inst_bytes	[736][0]	= 8'hD1;
		inst_bytes	[736][1]	= 8'hF9;
		inst_size	[736]		= 4'd2;

		inst_bytes	[737][0]	= 8'hD3;
		inst_bytes	[737][1]	= 8'h39;
		inst_size	[737]		= 4'd2;

		inst_bytes	[738][0]	= 8'hD3;
		inst_bytes	[738][1]	= 8'h3C;
		inst_bytes	[738][2]	= 8'h52;
		inst_size	[738]		= 4'd3;

		inst_bytes	[739][0]	= 8'hD3;
		inst_bytes	[739][1]	= 8'h3D;
		inst_bytes	[739][2]	= 8'h01;
		inst_bytes	[739][3]	= 8'h02;
		inst_bytes	[739][4]	= 8'h03;
		inst_bytes	[739][5]	= 8'h04;
		inst_size	[739]		= 4'd6;

		inst_bytes	[740][0]	= 8'hD3;
		inst_bytes	[740][1]	= 8'h79;
		inst_bytes	[740][2]	= 8'h01;
		inst_size	[740]		= 4'd3;

		inst_bytes	[741][0]	= 8'hD3;
		inst_bytes	[741][1]	= 8'h7C;
		inst_bytes	[741][2]	= 8'h52;
		inst_bytes	[741][3]	= 8'h01;
		inst_size	[741]		= 4'd4;

		inst_bytes	[742][0]	= 8'hD3;
		inst_bytes	[742][1]	= 8'hB9;
		inst_bytes	[742][2]	= 8'h01;
		inst_bytes	[742][3]	= 8'h02;
		inst_bytes	[742][4]	= 8'h03;
		inst_bytes	[742][5]	= 8'h04;
		inst_size	[742]		= 4'd6;

		inst_bytes	[743][0]	= 8'hD3;
		inst_bytes	[743][1]	= 8'hBC;
		inst_bytes	[743][2]	= 8'h52;
		inst_bytes	[743][3]	= 8'h01;
		inst_bytes	[743][4]	= 8'h02;
		inst_bytes	[743][5]	= 8'h03;
		inst_bytes	[743][6]	= 8'h04;
		inst_size	[743]		= 4'd7;

		inst_bytes	[744][0]	= 8'hD3;
		inst_bytes	[744][1]	= 8'hF9;
		inst_size	[744]		= 4'd2;

		inst_bytes	[745][0]	= 8'hC1;
		inst_bytes	[745][1]	= 8'h39;
		inst_bytes	[745][2]	= 8'h11;
		inst_size	[745]		= 4'd3;

		inst_bytes	[746][0]	= 8'hC1;
		inst_bytes	[746][1]	= 8'h3C;
		inst_bytes	[746][2]	= 8'h52;
		inst_bytes	[746][3]	= 8'h11;
		inst_size	[746]		= 4'd4;

		inst_bytes	[747][0]	= 8'hC1;
		inst_bytes	[747][1]	= 8'h3D;
		inst_bytes	[747][2]	= 8'h01;
		inst_bytes	[747][3]	= 8'h02;
		inst_bytes	[747][4]	= 8'h03;
		inst_bytes	[747][5]	= 8'h04;
		inst_bytes	[747][6]	= 8'h11;
		inst_size	[747]		= 4'd7;

		inst_bytes	[748][0]	= 8'hC1;
		inst_bytes	[748][1]	= 8'h79;
		inst_bytes	[748][2]	= 8'h01;
		inst_bytes	[748][3]	= 8'h11;
		inst_size	[748]		= 4'd4;

		inst_bytes	[749][0]	= 8'hC1;
		inst_bytes	[749][1]	= 8'h7C;
		inst_bytes	[749][2]	= 8'h52;
		inst_bytes	[749][3]	= 8'h01;
		inst_bytes	[749][4]	= 8'h11;
		inst_size	[749]		= 4'd5;

		inst_bytes	[750][0]	= 8'hC1;
		inst_bytes	[750][1]	= 8'hB9;
		inst_bytes	[750][2]	= 8'h01;
		inst_bytes	[750][3]	= 8'h02;
		inst_bytes	[750][4]	= 8'h03;
		inst_bytes	[750][5]	= 8'h04;
		inst_bytes	[750][6]	= 8'h11;
		inst_size	[750]		= 4'd7;

		inst_bytes	[751][0]	= 8'hC1;
		inst_bytes	[751][1]	= 8'hBC;
		inst_bytes	[751][2]	= 8'h52;
		inst_bytes	[751][3]	= 8'h01;
		inst_bytes	[751][4]	= 8'h02;
		inst_bytes	[751][5]	= 8'h03;
		inst_bytes	[751][6]	= 8'h04;
		inst_bytes	[751][7]	= 8'h11;
		inst_size	[751]		= 4'd8;

		inst_bytes	[752][0]	= 8'hC1;
		inst_bytes	[752][1]	= 8'hF9;
		inst_bytes	[752][2]	= 8'h11;
		inst_size	[752]		= 4'd3;

		inst_bytes	[753][0]	= 8'hFD;
		inst_size	[753]		= 4'd1;

		inst_bytes	[754][0]	= 8'h66;
		inst_bytes	[754][1]	= 8'h91;
		inst_size	[754]		= 4'd2;

		inst_bytes	[755][0]	= 8'h91;
		inst_size	[755]		= 4'd1;

		inst_bytes	[756][0]	= 8'h86;
		inst_bytes	[756][1]	= 8'h01;
		inst_size	[756]		= 4'd2;

		inst_bytes	[757][0]	= 8'h86;
		inst_bytes	[757][1]	= 8'h04;
		inst_bytes	[757][2]	= 8'h52;
		inst_size	[757]		= 4'd3;

		inst_bytes	[758][0]	= 8'h86;
		inst_bytes	[758][1]	= 8'h05;
		inst_bytes	[758][2]	= 8'h01;
		inst_bytes	[758][3]	= 8'h02;
		inst_bytes	[758][4]	= 8'h03;
		inst_bytes	[758][5]	= 8'h04;
		inst_size	[758]		= 4'd6;

		inst_bytes	[759][0]	= 8'h86;
		inst_bytes	[759][1]	= 8'h41;
		inst_bytes	[759][2]	= 8'h01;
		inst_size	[759]		= 4'd3;

		inst_bytes	[760][0]	= 8'h86;
		inst_bytes	[760][1]	= 8'h44;
		inst_bytes	[760][2]	= 8'h52;
		inst_bytes	[760][3]	= 8'h01;
		inst_size	[760]		= 4'd4;

		inst_bytes	[761][0]	= 8'h86;
		inst_bytes	[761][1]	= 8'h81;
		inst_bytes	[761][2]	= 8'h01;
		inst_bytes	[761][3]	= 8'h02;
		inst_bytes	[761][4]	= 8'h03;
		inst_bytes	[761][5]	= 8'h04;
		inst_size	[761]		= 4'd6;

		inst_bytes	[762][0]	= 8'h86;
		inst_bytes	[762][1]	= 8'h84;
		inst_bytes	[762][2]	= 8'h52;
		inst_bytes	[762][3]	= 8'h01;
		inst_bytes	[762][4]	= 8'h02;
		inst_bytes	[762][5]	= 8'h03;
		inst_bytes	[762][6]	= 8'h04;
		inst_size	[762]		= 4'd7;

		inst_bytes	[763][0]	= 8'h86;
		inst_bytes	[763][1]	= 8'hC1;
		inst_size	[763]		= 4'd2;

		inst_bytes	[764][0]	= 8'h87;
		inst_bytes	[764][1]	= 8'h01;
		inst_size	[764]		= 4'd2;

		inst_bytes	[765][0]	= 8'h87;
		inst_bytes	[765][1]	= 8'h04;
		inst_bytes	[765][2]	= 8'h52;
		inst_size	[765]		= 4'd3;

		inst_bytes	[766][0]	= 8'h87;
		inst_bytes	[766][1]	= 8'h05;
		inst_bytes	[766][2]	= 8'h01;
		inst_bytes	[766][3]	= 8'h02;
		inst_bytes	[766][4]	= 8'h03;
		inst_bytes	[766][5]	= 8'h04;
		inst_size	[766]		= 4'd6;

		inst_bytes	[767][0]	= 8'h87;
		inst_bytes	[767][1]	= 8'h41;
		inst_bytes	[767][2]	= 8'h01;
		inst_size	[767]		= 4'd3;

		inst_bytes	[768][0]	= 8'h87;
		inst_bytes	[768][1]	= 8'h44;
		inst_bytes	[768][2]	= 8'h52;
		inst_bytes	[768][3]	= 8'h01;
		inst_size	[768]		= 4'd4;

		inst_bytes	[769][0]	= 8'h87;
		inst_bytes	[769][1]	= 8'h81;
		inst_bytes	[769][2]	= 8'h01;
		inst_bytes	[769][3]	= 8'h02;
		inst_bytes	[769][4]	= 8'h03;
		inst_bytes	[769][5]	= 8'h04;
		inst_size	[769]		= 4'd6;

		inst_bytes	[770][0]	= 8'h87;
		inst_bytes	[770][1]	= 8'h84;
		inst_bytes	[770][2]	= 8'h52;
		inst_bytes	[770][3]	= 8'h01;
		inst_bytes	[770][4]	= 8'h02;
		inst_bytes	[770][5]	= 8'h03;
		inst_bytes	[770][6]	= 8'h04;
		inst_size	[770]		= 4'd7;

		inst_bytes	[771][0]	= 8'h87;
		inst_bytes	[771][1]	= 8'hC1;
		inst_size	[771]		= 4'd2;

		inst_bytes	[772][0]	= 8'h87;
		inst_bytes	[772][1]	= 8'h01;
		inst_size	[772]		= 4'd2;

		inst_bytes	[773][0]	= 8'h87;
		inst_bytes	[773][1]	= 8'h04;
		inst_bytes	[773][2]	= 8'h52;
		inst_size	[773]		= 4'd3;

		inst_bytes	[774][0]	= 8'h87;
		inst_bytes	[774][1]	= 8'h05;
		inst_bytes	[774][2]	= 8'h01;
		inst_bytes	[774][3]	= 8'h02;
		inst_bytes	[774][4]	= 8'h03;
		inst_bytes	[774][5]	= 8'h04;
		inst_size	[774]		= 4'd6;

		inst_bytes	[775][0]	= 8'h87;
		inst_bytes	[775][1]	= 8'h41;
		inst_bytes	[775][2]	= 8'h01;
		inst_size	[775]		= 4'd3;

		inst_bytes	[776][0]	= 8'h87;
		inst_bytes	[776][1]	= 8'h44;
		inst_bytes	[776][2]	= 8'h52;
		inst_bytes	[776][3]	= 8'h01;
		inst_size	[776]		= 4'd4;

		inst_bytes	[777][0]	= 8'h87;
		inst_bytes	[777][1]	= 8'h81;
		inst_bytes	[777][2]	= 8'h01;
		inst_bytes	[777][3]	= 8'h02;
		inst_bytes	[777][4]	= 8'h03;
		inst_bytes	[777][5]	= 8'h04;
		inst_size	[777]		= 4'd6;

		inst_bytes	[778][0]	= 8'h87;
		inst_bytes	[778][1]	= 8'h84;
		inst_bytes	[778][2]	= 8'h52;
		inst_bytes	[778][3]	= 8'h01;
		inst_bytes	[778][4]	= 8'h02;
		inst_bytes	[778][5]	= 8'h03;
		inst_bytes	[778][6]	= 8'h04;
		inst_size	[778]		= 4'd7;

		inst_bytes	[779][0]	= 8'h87;
		inst_bytes	[779][1]	= 8'hC1;
		inst_size	[779]		= 4'd2;

	end


	reg	[63:0]	cache_lines	[447:0];
	initial begin

		cache_lines[0]		= {inst_bytes[0][0], inst_bytes[0][1], inst_bytes[1][0], inst_bytes[1][1], inst_bytes[1][2], inst_bytes[1][3], inst_bytes[2][0], inst_bytes[2][1]};

		cache_lines[1]		= {inst_bytes[2][2], inst_bytes[2][3], inst_bytes[2][4], inst_bytes[3][0], inst_bytes[3][1], inst_bytes[3][2], inst_bytes[4][0], inst_bytes[4][1]};

		cache_lines[2]		= {inst_bytes[4][2], inst_bytes[4][3], inst_bytes[5][0], inst_bytes[5][1], inst_bytes[5][2], inst_bytes[5][3], inst_bytes[5][4], inst_bytes[5][5]};

		cache_lines[3]		= {inst_bytes[5][6], inst_bytes[6][0], inst_bytes[6][1], inst_bytes[6][2], inst_bytes[6][3], inst_bytes[7][0], inst_bytes[7][1], inst_bytes[7][2]};

		cache_lines[4]		= {inst_bytes[7][3], inst_bytes[7][4], inst_bytes[8][0], inst_bytes[8][1], inst_bytes[8][2], inst_bytes[8][3], inst_bytes[8][4], inst_bytes[8][5]};

		cache_lines[5]		= {inst_bytes[8][6], inst_bytes[9][0], inst_bytes[9][1], inst_bytes[9][2], inst_bytes[9][3], inst_bytes[9][4], inst_bytes[9][5], inst_bytes[9][6]};

		cache_lines[6]		= {inst_bytes[9][7], inst_bytes[10][0], inst_bytes[10][1], inst_bytes[10][2], inst_bytes[11][0], inst_bytes[11][1], inst_bytes[11][2], inst_bytes[11][3]};

		cache_lines[7]		= {inst_bytes[11][4], inst_bytes[12][0], inst_bytes[12][1], inst_bytes[12][2], inst_bytes[12][3], inst_bytes[12][4], inst_bytes[12][5], inst_bytes[13][0]};

		cache_lines[8]		= {inst_bytes[13][1], inst_bytes[13][2], inst_bytes[13][3], inst_bytes[13][4], inst_bytes[13][5], inst_bytes[13][6], inst_bytes[13][7], inst_bytes[13][8]};

		cache_lines[9]		= {inst_bytes[14][0], inst_bytes[14][1], inst_bytes[14][2], inst_bytes[14][3], inst_bytes[14][4], inst_bytes[14][5], inst_bytes[15][0], inst_bytes[15][1]};

		cache_lines[10]		= {inst_bytes[15][2], inst_bytes[15][3], inst_bytes[15][4], inst_bytes[15][5], inst_bytes[15][6], inst_bytes[16][0], inst_bytes[16][1], inst_bytes[16][2]};

		cache_lines[11]		= {inst_bytes[16][3], inst_bytes[16][4], inst_bytes[16][5], inst_bytes[16][6], inst_bytes[16][7], inst_bytes[16][8], inst_bytes[17][0], inst_bytes[17][1]};

		cache_lines[12]		= {inst_bytes[17][2], inst_bytes[17][3], inst_bytes[17][4], inst_bytes[17][5], inst_bytes[17][6], inst_bytes[17][7], inst_bytes[17][8], inst_bytes[17][9]};

		cache_lines[13]		= {inst_bytes[18][0], inst_bytes[18][1], inst_bytes[18][2], inst_bytes[18][3], inst_bytes[18][4], inst_bytes[19][0], inst_bytes[19][1], inst_bytes[19][2]};

		cache_lines[14]		= {inst_bytes[19][3], inst_bytes[19][4], inst_bytes[19][5], inst_bytes[20][0], inst_bytes[20][1], inst_bytes[20][2], inst_bytes[20][3], inst_bytes[20][4]};

		cache_lines[15]		= {inst_bytes[20][5], inst_bytes[20][6], inst_bytes[21][0], inst_bytes[21][1], inst_bytes[21][2], inst_bytes[21][3], inst_bytes[21][4], inst_bytes[21][5]};

		cache_lines[16]		= {inst_bytes[21][6], inst_bytes[21][7], inst_bytes[21][8], inst_bytes[21][9], inst_bytes[22][0], inst_bytes[22][1], inst_bytes[22][2], inst_bytes[22][3]};

		cache_lines[17]		= {inst_bytes[22][4], inst_bytes[22][5], inst_bytes[22][6], inst_bytes[23][0], inst_bytes[23][1], inst_bytes[23][2], inst_bytes[23][3], inst_bytes[23][4]};

		cache_lines[18]		= {inst_bytes[23][5], inst_bytes[23][6], inst_bytes[23][7], inst_bytes[24][0], inst_bytes[24][1], inst_bytes[24][2], inst_bytes[24][3], inst_bytes[24][4]};

		cache_lines[19]		= {inst_bytes[24][5], inst_bytes[24][6], inst_bytes[24][7], inst_bytes[24][8], inst_bytes[24][9], inst_bytes[25][0], inst_bytes[25][1], inst_bytes[25][2]};

		cache_lines[20]		= {inst_bytes[25][3], inst_bytes[25][4], inst_bytes[25][5], inst_bytes[25][6], inst_bytes[25][7], inst_bytes[25][8], inst_bytes[25][9], inst_bytes[25][10]};

		cache_lines[21]		= {inst_bytes[26][0], inst_bytes[26][1], inst_bytes[26][2], inst_bytes[26][3], inst_bytes[26][4], inst_bytes[26][5], inst_bytes[27][0], inst_bytes[27][1]};

		cache_lines[22]		= {inst_bytes[27][2], inst_bytes[28][0], inst_bytes[28][1], inst_bytes[28][2], inst_bytes[28][3], inst_bytes[29][0], inst_bytes[29][1], inst_bytes[29][2]};

		cache_lines[23]		= {inst_bytes[29][3], inst_bytes[29][4], inst_bytes[29][5], inst_bytes[29][6], inst_bytes[30][0], inst_bytes[30][1], inst_bytes[30][2], inst_bytes[30][3]};

		cache_lines[24]		= {inst_bytes[31][0], inst_bytes[31][1], inst_bytes[31][2], inst_bytes[31][3], inst_bytes[31][4], inst_bytes[32][0], inst_bytes[32][1], inst_bytes[32][2]};

		cache_lines[25]		= {inst_bytes[32][3], inst_bytes[32][4], inst_bytes[32][5], inst_bytes[32][6], inst_bytes[33][0], inst_bytes[33][1], inst_bytes[33][2], inst_bytes[33][3]};

		cache_lines[26]		= {inst_bytes[33][4], inst_bytes[33][5], inst_bytes[33][6], inst_bytes[33][7], inst_bytes[34][0], inst_bytes[34][1], inst_bytes[34][2], inst_bytes[35][0]};

		cache_lines[27]		= {inst_bytes[35][1], inst_bytes[35][2], inst_bytes[36][0], inst_bytes[36][1], inst_bytes[36][2], inst_bytes[36][3], inst_bytes[37][0], inst_bytes[37][1]};

		cache_lines[28]		= {inst_bytes[37][2], inst_bytes[37][3], inst_bytes[37][4], inst_bytes[37][5], inst_bytes[37][6], inst_bytes[38][0], inst_bytes[38][1], inst_bytes[38][2]};

		cache_lines[29]		= {inst_bytes[38][3], inst_bytes[39][0], inst_bytes[39][1], inst_bytes[39][2], inst_bytes[39][3], inst_bytes[39][4], inst_bytes[40][0], inst_bytes[40][1]};

		cache_lines[30]		= {inst_bytes[40][2], inst_bytes[40][3], inst_bytes[40][4], inst_bytes[40][5], inst_bytes[40][6], inst_bytes[41][0], inst_bytes[41][1], inst_bytes[41][2]};

		cache_lines[31]		= {inst_bytes[41][3], inst_bytes[41][4], inst_bytes[41][5], inst_bytes[41][6], inst_bytes[41][7], inst_bytes[42][0], inst_bytes[42][1], inst_bytes[42][2]};

		cache_lines[32]		= {inst_bytes[43][0], inst_bytes[43][1], inst_bytes[44][0], inst_bytes[44][1], inst_bytes[44][2], inst_bytes[45][0], inst_bytes[45][1], inst_bytes[45][2]};

		cache_lines[33]		= {inst_bytes[45][3], inst_bytes[45][4], inst_bytes[45][5], inst_bytes[46][0], inst_bytes[46][1], inst_bytes[46][2], inst_bytes[47][0], inst_bytes[47][1]};

		cache_lines[34]		= {inst_bytes[47][2], inst_bytes[47][3], inst_bytes[48][0], inst_bytes[48][1], inst_bytes[48][2], inst_bytes[48][3], inst_bytes[48][4], inst_bytes[48][5]};

		cache_lines[35]		= {inst_bytes[49][0], inst_bytes[49][1], inst_bytes[49][2], inst_bytes[49][3], inst_bytes[49][4], inst_bytes[49][5], inst_bytes[49][6], inst_bytes[50][0]};

		cache_lines[36]		= {inst_bytes[50][1], inst_bytes[51][0], inst_bytes[51][1], inst_bytes[52][0], inst_bytes[52][1], inst_bytes[52][2], inst_bytes[53][0], inst_bytes[53][1]};

		cache_lines[37]		= {inst_bytes[53][2], inst_bytes[53][3], inst_bytes[53][4], inst_bytes[53][5], inst_bytes[54][0], inst_bytes[54][1], inst_bytes[54][2], inst_bytes[55][0]};

		cache_lines[38]		= {inst_bytes[55][1], inst_bytes[55][2], inst_bytes[55][3], inst_bytes[56][0], inst_bytes[56][1], inst_bytes[56][2], inst_bytes[56][3], inst_bytes[56][4]};

		cache_lines[39]		= {inst_bytes[56][5], inst_bytes[57][0], inst_bytes[57][1], inst_bytes[57][2], inst_bytes[57][3], inst_bytes[57][4], inst_bytes[57][5], inst_bytes[57][6]};

		cache_lines[40]		= {inst_bytes[58][0], inst_bytes[58][1], inst_bytes[59][0], inst_bytes[59][1], inst_bytes[60][0], inst_bytes[60][1], inst_bytes[60][2], inst_bytes[61][0]};

		cache_lines[41]		= {inst_bytes[61][1], inst_bytes[61][2], inst_bytes[61][3], inst_bytes[61][4], inst_bytes[61][5], inst_bytes[62][0], inst_bytes[62][1], inst_bytes[62][2]};

		cache_lines[42]		= {inst_bytes[63][0], inst_bytes[63][1], inst_bytes[63][2], inst_bytes[63][3], inst_bytes[64][0], inst_bytes[64][1], inst_bytes[64][2], inst_bytes[64][3]};

		cache_lines[43]		= {inst_bytes[64][4], inst_bytes[64][5], inst_bytes[65][0], inst_bytes[65][1], inst_bytes[65][2], inst_bytes[65][3], inst_bytes[65][4], inst_bytes[65][5]};

		cache_lines[44]		= {inst_bytes[65][6], inst_bytes[66][0], inst_bytes[66][1], inst_bytes[67][0], inst_bytes[67][1], inst_bytes[68][0], inst_bytes[68][1], inst_bytes[68][2]};

		cache_lines[45]		= {inst_bytes[69][0], inst_bytes[69][1], inst_bytes[69][2], inst_bytes[69][3], inst_bytes[69][4], inst_bytes[69][5], inst_bytes[70][0], inst_bytes[70][1]};

		cache_lines[46]		= {inst_bytes[70][2], inst_bytes[71][0], inst_bytes[71][1], inst_bytes[71][2], inst_bytes[71][3], inst_bytes[72][0], inst_bytes[72][1], inst_bytes[72][2]};

		cache_lines[47]		= {inst_bytes[72][3], inst_bytes[72][4], inst_bytes[72][5], inst_bytes[73][0], inst_bytes[73][1], inst_bytes[73][2], inst_bytes[73][3], inst_bytes[73][4]};

		cache_lines[48]		= {inst_bytes[73][5], inst_bytes[73][6], inst_bytes[74][0], inst_bytes[74][1], inst_bytes[75][0], inst_bytes[75][1], inst_bytes[76][0], inst_bytes[76][1]};

		cache_lines[49]		= {inst_bytes[76][2], inst_bytes[77][0], inst_bytes[77][1], inst_bytes[77][2], inst_bytes[77][3], inst_bytes[77][4], inst_bytes[77][5], inst_bytes[78][0]};

		cache_lines[50]		= {inst_bytes[78][1], inst_bytes[78][2], inst_bytes[79][0], inst_bytes[79][1], inst_bytes[79][2], inst_bytes[79][3], inst_bytes[80][0], inst_bytes[80][1]};

		cache_lines[51]		= {inst_bytes[80][2], inst_bytes[80][3], inst_bytes[80][4], inst_bytes[80][5], inst_bytes[81][0], inst_bytes[81][1], inst_bytes[81][2], inst_bytes[81][3]};

		cache_lines[52]		= {inst_bytes[81][4], inst_bytes[81][5], inst_bytes[81][6], inst_bytes[82][0], inst_bytes[82][1], inst_bytes[83][0], inst_bytes[83][1], inst_bytes[84][0]};

		cache_lines[53]		= {inst_bytes[84][1], inst_bytes[84][2], inst_bytes[85][0], inst_bytes[85][1], inst_bytes[85][2], inst_bytes[85][3], inst_bytes[85][4], inst_bytes[85][5]};

		cache_lines[54]		= {inst_bytes[86][0], inst_bytes[86][1], inst_bytes[86][2], inst_bytes[87][0], inst_bytes[87][1], inst_bytes[87][2], inst_bytes[87][3], inst_bytes[88][0]};

		cache_lines[55]		= {inst_bytes[88][1], inst_bytes[88][2], inst_bytes[88][3], inst_bytes[88][4], inst_bytes[88][5], inst_bytes[89][0], inst_bytes[89][1], inst_bytes[89][2]};

		cache_lines[56]		= {inst_bytes[89][3], inst_bytes[89][4], inst_bytes[89][5], inst_bytes[89][6], inst_bytes[90][0], inst_bytes[90][1], inst_bytes[91][0], inst_bytes[91][1]};

		cache_lines[57]		= {inst_bytes[92][0], inst_bytes[92][1], inst_bytes[92][2], inst_bytes[92][3], inst_bytes[93][0], inst_bytes[93][1], inst_bytes[93][2], inst_bytes[93][3]};

		cache_lines[58]		= {inst_bytes[93][4], inst_bytes[94][0], inst_bytes[94][1], inst_bytes[94][2], inst_bytes[95][0], inst_bytes[95][1], inst_bytes[95][2], inst_bytes[95][3]};

		cache_lines[59]		= {inst_bytes[96][0], inst_bytes[96][1], inst_bytes[96][2], inst_bytes[96][3], inst_bytes[96][4], inst_bytes[96][5], inst_bytes[96][6], inst_bytes[97][0]};

		cache_lines[60]		= {inst_bytes[97][1], inst_bytes[97][2], inst_bytes[97][3], inst_bytes[98][0], inst_bytes[98][1], inst_bytes[98][2], inst_bytes[98][3], inst_bytes[98][4]};

		cache_lines[61]		= {inst_bytes[99][0], inst_bytes[99][1], inst_bytes[99][2], inst_bytes[99][3], inst_bytes[99][4], inst_bytes[99][5], inst_bytes[99][6], inst_bytes[100][0]};

		cache_lines[62]		= {inst_bytes[100][1], inst_bytes[100][2], inst_bytes[100][3], inst_bytes[100][4], inst_bytes[100][5], inst_bytes[100][6], inst_bytes[100][7], inst_bytes[101][0]};

		cache_lines[63]		= {inst_bytes[101][1], inst_bytes[101][2], inst_bytes[102][0], inst_bytes[102][1], inst_bytes[102][2], inst_bytes[102][3], inst_bytes[102][4], inst_bytes[103][0]};

		cache_lines[64]		= {inst_bytes[103][1], inst_bytes[103][2], inst_bytes[103][3], inst_bytes[103][4], inst_bytes[103][5], inst_bytes[104][0], inst_bytes[104][1], inst_bytes[104][2]};

		cache_lines[65]		= {inst_bytes[104][3], inst_bytes[104][4], inst_bytes[104][5], inst_bytes[104][6], inst_bytes[104][7], inst_bytes[104][8], inst_bytes[105][0], inst_bytes[105][1]};

		cache_lines[66]		= {inst_bytes[105][2], inst_bytes[105][3], inst_bytes[105][4], inst_bytes[105][5], inst_bytes[106][0], inst_bytes[106][1], inst_bytes[106][2], inst_bytes[106][3]};

		cache_lines[67]		= {inst_bytes[106][4], inst_bytes[106][5], inst_bytes[106][6], inst_bytes[107][0], inst_bytes[107][1], inst_bytes[107][2], inst_bytes[107][3], inst_bytes[107][4]};

		cache_lines[68]		= {inst_bytes[107][5], inst_bytes[107][6], inst_bytes[107][7], inst_bytes[107][8], inst_bytes[108][0], inst_bytes[108][1], inst_bytes[108][2], inst_bytes[108][3]};

		cache_lines[69]		= {inst_bytes[108][4], inst_bytes[108][5], inst_bytes[108][6], inst_bytes[108][7], inst_bytes[108][8], inst_bytes[108][9], inst_bytes[109][0], inst_bytes[109][1]};

		cache_lines[70]		= {inst_bytes[109][2], inst_bytes[109][3], inst_bytes[109][4], inst_bytes[110][0], inst_bytes[110][1], inst_bytes[110][2], inst_bytes[110][3], inst_bytes[110][4]};

		cache_lines[71]		= {inst_bytes[110][5], inst_bytes[111][0], inst_bytes[111][1], inst_bytes[111][2], inst_bytes[111][3], inst_bytes[111][4], inst_bytes[111][5], inst_bytes[111][6]};

		cache_lines[72]		= {inst_bytes[112][0], inst_bytes[112][1], inst_bytes[112][2], inst_bytes[112][3], inst_bytes[112][4], inst_bytes[112][5], inst_bytes[112][6], inst_bytes[112][7]};

		cache_lines[73]		= {inst_bytes[112][8], inst_bytes[112][9], inst_bytes[113][0], inst_bytes[113][1], inst_bytes[113][2], inst_bytes[113][3], inst_bytes[113][4], inst_bytes[113][5]};

		cache_lines[74]		= {inst_bytes[113][6], inst_bytes[114][0], inst_bytes[114][1], inst_bytes[114][2], inst_bytes[114][3], inst_bytes[114][4], inst_bytes[114][5], inst_bytes[114][6]};

		cache_lines[75]		= {inst_bytes[114][7], inst_bytes[115][0], inst_bytes[115][1], inst_bytes[115][2], inst_bytes[115][3], inst_bytes[115][4], inst_bytes[115][5], inst_bytes[115][6]};

		cache_lines[76]		= {inst_bytes[115][7], inst_bytes[115][8], inst_bytes[115][9], inst_bytes[116][0], inst_bytes[116][1], inst_bytes[116][2], inst_bytes[116][3], inst_bytes[116][4]};

		cache_lines[77]		= {inst_bytes[116][5], inst_bytes[116][6], inst_bytes[116][7], inst_bytes[116][8], inst_bytes[116][9], inst_bytes[116][10], inst_bytes[117][0], inst_bytes[117][1]};

		cache_lines[78]		= {inst_bytes[117][2], inst_bytes[117][3], inst_bytes[117][4], inst_bytes[117][5], inst_bytes[118][0], inst_bytes[118][1], inst_bytes[118][2], inst_bytes[119][0]};

		cache_lines[79]		= {inst_bytes[119][1], inst_bytes[119][2], inst_bytes[119][3], inst_bytes[120][0], inst_bytes[120][1], inst_bytes[120][2], inst_bytes[120][3], inst_bytes[120][4]};

		cache_lines[80]		= {inst_bytes[120][5], inst_bytes[120][6], inst_bytes[121][0], inst_bytes[121][1], inst_bytes[121][2], inst_bytes[121][3], inst_bytes[122][0], inst_bytes[122][1]};

		cache_lines[81]		= {inst_bytes[122][2], inst_bytes[122][3], inst_bytes[122][4], inst_bytes[123][0], inst_bytes[123][1], inst_bytes[123][2], inst_bytes[123][3], inst_bytes[123][4]};

		cache_lines[82]		= {inst_bytes[123][5], inst_bytes[123][6], inst_bytes[124][0], inst_bytes[124][1], inst_bytes[124][2], inst_bytes[124][3], inst_bytes[124][4], inst_bytes[124][5]};

		cache_lines[83]		= {inst_bytes[124][6], inst_bytes[124][7], inst_bytes[125][0], inst_bytes[125][1], inst_bytes[125][2], inst_bytes[126][0], inst_bytes[126][1], inst_bytes[126][2]};

		cache_lines[84]		= {inst_bytes[127][0], inst_bytes[127][1], inst_bytes[127][2], inst_bytes[127][3], inst_bytes[128][0], inst_bytes[128][1], inst_bytes[128][2], inst_bytes[128][3]};

		cache_lines[85]		= {inst_bytes[128][4], inst_bytes[128][5], inst_bytes[128][6], inst_bytes[129][0], inst_bytes[129][1], inst_bytes[129][2], inst_bytes[129][3], inst_bytes[130][0]};

		cache_lines[86]		= {inst_bytes[130][1], inst_bytes[130][2], inst_bytes[130][3], inst_bytes[130][4], inst_bytes[131][0], inst_bytes[131][1], inst_bytes[131][2], inst_bytes[131][3]};

		cache_lines[87]		= {inst_bytes[131][4], inst_bytes[131][5], inst_bytes[131][6], inst_bytes[132][0], inst_bytes[132][1], inst_bytes[132][2], inst_bytes[132][3], inst_bytes[132][4]};

		cache_lines[88]		= {inst_bytes[132][5], inst_bytes[132][6], inst_bytes[132][7], inst_bytes[133][0], inst_bytes[133][1], inst_bytes[133][2], inst_bytes[134][0], inst_bytes[134][1]};

		cache_lines[89]		= {inst_bytes[135][0], inst_bytes[135][1], inst_bytes[135][2], inst_bytes[136][0], inst_bytes[136][1], inst_bytes[136][2], inst_bytes[136][3], inst_bytes[136][4]};

		cache_lines[90]		= {inst_bytes[136][5], inst_bytes[137][0], inst_bytes[137][1], inst_bytes[137][2], inst_bytes[138][0], inst_bytes[138][1], inst_bytes[138][2], inst_bytes[138][3]};

		cache_lines[91]		= {inst_bytes[139][0], inst_bytes[139][1], inst_bytes[139][2], inst_bytes[139][3], inst_bytes[139][4], inst_bytes[139][5], inst_bytes[140][0], inst_bytes[140][1]};

		cache_lines[92]		= {inst_bytes[140][2], inst_bytes[140][3], inst_bytes[140][4], inst_bytes[140][5], inst_bytes[140][6], inst_bytes[141][0], inst_bytes[141][1], inst_bytes[142][0]};

		cache_lines[93]		= {inst_bytes[142][1], inst_bytes[143][0], inst_bytes[143][1], inst_bytes[143][2], inst_bytes[144][0], inst_bytes[144][1], inst_bytes[144][2], inst_bytes[144][3]};

		cache_lines[94]		= {inst_bytes[144][4], inst_bytes[144][5], inst_bytes[145][0], inst_bytes[145][1], inst_bytes[145][2], inst_bytes[146][0], inst_bytes[146][1], inst_bytes[146][2]};

		cache_lines[95]		= {inst_bytes[146][3], inst_bytes[147][0], inst_bytes[147][1], inst_bytes[147][2], inst_bytes[147][3], inst_bytes[147][4], inst_bytes[147][5], inst_bytes[148][0]};

		cache_lines[96]		= {inst_bytes[148][1], inst_bytes[148][2], inst_bytes[148][3], inst_bytes[148][4], inst_bytes[148][5], inst_bytes[148][6], inst_bytes[149][0], inst_bytes[149][1]};

		cache_lines[97]		= {inst_bytes[150][0], inst_bytes[150][1], inst_bytes[151][0], inst_bytes[151][1], inst_bytes[151][2], inst_bytes[152][0], inst_bytes[152][1], inst_bytes[152][2]};

		cache_lines[98]		= {inst_bytes[152][3], inst_bytes[152][4], inst_bytes[152][5], inst_bytes[153][0], inst_bytes[153][1], inst_bytes[153][2], inst_bytes[154][0], inst_bytes[154][1]};

		cache_lines[99]		= {inst_bytes[154][2], inst_bytes[154][3], inst_bytes[155][0], inst_bytes[155][1], inst_bytes[155][2], inst_bytes[155][3], inst_bytes[155][4], inst_bytes[155][5]};

		cache_lines[100]		= {inst_bytes[156][0], inst_bytes[156][1], inst_bytes[156][2], inst_bytes[156][3], inst_bytes[156][4], inst_bytes[156][5], inst_bytes[156][6], inst_bytes[157][0]};

		cache_lines[101]		= {inst_bytes[157][1], inst_bytes[158][0], inst_bytes[158][1], inst_bytes[159][0], inst_bytes[159][1], inst_bytes[159][2], inst_bytes[160][0], inst_bytes[160][1]};

		cache_lines[102]		= {inst_bytes[160][2], inst_bytes[160][3], inst_bytes[160][4], inst_bytes[160][5], inst_bytes[161][0], inst_bytes[161][1], inst_bytes[161][2], inst_bytes[162][0]};

		cache_lines[103]		= {inst_bytes[162][1], inst_bytes[162][2], inst_bytes[162][3], inst_bytes[163][0], inst_bytes[163][1], inst_bytes[163][2], inst_bytes[163][3], inst_bytes[163][4]};

		cache_lines[104]		= {inst_bytes[163][5], inst_bytes[164][0], inst_bytes[164][1], inst_bytes[164][2], inst_bytes[164][3], inst_bytes[164][4], inst_bytes[164][5], inst_bytes[164][6]};

		cache_lines[105]		= {inst_bytes[165][0], inst_bytes[165][1], inst_bytes[166][0], inst_bytes[166][1], inst_bytes[167][0], inst_bytes[167][1], inst_bytes[167][2], inst_bytes[168][0]};

		cache_lines[106]		= {inst_bytes[168][1], inst_bytes[168][2], inst_bytes[168][3], inst_bytes[168][4], inst_bytes[168][5], inst_bytes[169][0], inst_bytes[169][1], inst_bytes[169][2]};

		cache_lines[107]		= {inst_bytes[170][0], inst_bytes[170][1], inst_bytes[170][2], inst_bytes[170][3], inst_bytes[171][0], inst_bytes[171][1], inst_bytes[171][2], inst_bytes[171][3]};

		cache_lines[108]		= {inst_bytes[171][4], inst_bytes[171][5], inst_bytes[172][0], inst_bytes[172][1], inst_bytes[172][2], inst_bytes[172][3], inst_bytes[172][4], inst_bytes[172][5]};

		cache_lines[109]		= {inst_bytes[172][6], inst_bytes[173][0], inst_bytes[173][1], inst_bytes[174][0], inst_bytes[174][1], inst_bytes[175][0], inst_bytes[175][1], inst_bytes[175][2]};

		cache_lines[110]		= {inst_bytes[176][0], inst_bytes[176][1], inst_bytes[176][2], inst_bytes[176][3], inst_bytes[176][4], inst_bytes[176][5], inst_bytes[177][0], inst_bytes[177][1]};

		cache_lines[111]		= {inst_bytes[177][2], inst_bytes[178][0], inst_bytes[178][1], inst_bytes[178][2], inst_bytes[178][3], inst_bytes[179][0], inst_bytes[179][1], inst_bytes[179][2]};

		cache_lines[112]		= {inst_bytes[179][3], inst_bytes[179][4], inst_bytes[179][5], inst_bytes[180][0], inst_bytes[180][1], inst_bytes[180][2], inst_bytes[180][3], inst_bytes[180][4]};

		cache_lines[113]		= {inst_bytes[180][5], inst_bytes[180][6], inst_bytes[181][0], inst_bytes[181][1], inst_bytes[182][0], inst_bytes[182][1], inst_bytes[182][2], inst_bytes[182][3]};

		cache_lines[114]		= {inst_bytes[183][0], inst_bytes[183][1], inst_bytes[183][2], inst_bytes[183][3], inst_bytes[183][4], inst_bytes[184][0], inst_bytes[184][1], inst_bytes[185][0]};

		cache_lines[115]		= {inst_bytes[185][1], inst_bytes[185][2], inst_bytes[186][0], inst_bytes[186][1], inst_bytes[186][2], inst_bytes[186][3], inst_bytes[186][4], inst_bytes[186][5]};

		cache_lines[116]		= {inst_bytes[187][0], inst_bytes[187][1], inst_bytes[187][2], inst_bytes[188][0], inst_bytes[188][1], inst_bytes[188][2], inst_bytes[188][3], inst_bytes[189][0]};

		cache_lines[117]		= {inst_bytes[189][1], inst_bytes[189][2], inst_bytes[189][3], inst_bytes[189][4], inst_bytes[189][5], inst_bytes[190][0], inst_bytes[190][1], inst_bytes[190][2]};

		cache_lines[118]		= {inst_bytes[190][3], inst_bytes[190][4], inst_bytes[190][5], inst_bytes[190][6], inst_bytes[191][0], inst_bytes[191][1], inst_bytes[192][0], inst_bytes[192][1]};

		cache_lines[119]		= {inst_bytes[193][0], inst_bytes[193][1], inst_bytes[193][2], inst_bytes[194][0], inst_bytes[194][1], inst_bytes[194][2], inst_bytes[194][3], inst_bytes[194][4]};

		cache_lines[120]		= {inst_bytes[194][5], inst_bytes[195][0], inst_bytes[195][1], inst_bytes[195][2], inst_bytes[196][0], inst_bytes[196][1], inst_bytes[196][2], inst_bytes[196][3]};

		cache_lines[121]		= {inst_bytes[197][0], inst_bytes[197][1], inst_bytes[197][2], inst_bytes[197][3], inst_bytes[197][4], inst_bytes[197][5], inst_bytes[198][0], inst_bytes[198][1]};

		cache_lines[122]		= {inst_bytes[198][2], inst_bytes[198][3], inst_bytes[198][4], inst_bytes[198][5], inst_bytes[198][6], inst_bytes[199][0], inst_bytes[199][1], inst_bytes[200][0]};

		cache_lines[123]		= {inst_bytes[200][1], inst_bytes[200][2], inst_bytes[200][3], inst_bytes[200][4], inst_bytes[200][5], inst_bytes[200][6], inst_bytes[201][0], inst_bytes[202][0]};

		cache_lines[124]		= {inst_bytes[202][1], inst_bytes[202][2], inst_bytes[203][0], inst_bytes[203][1], inst_bytes[203][2], inst_bytes[203][3], inst_bytes[204][0], inst_bytes[204][1]};

		cache_lines[125]		= {inst_bytes[204][2], inst_bytes[204][3], inst_bytes[204][4], inst_bytes[204][5], inst_bytes[204][6], inst_bytes[205][0], inst_bytes[205][1], inst_bytes[205][2]};

		cache_lines[126]		= {inst_bytes[205][3], inst_bytes[206][0], inst_bytes[206][1], inst_bytes[206][2], inst_bytes[206][3], inst_bytes[206][4], inst_bytes[207][0], inst_bytes[207][1]};

		cache_lines[127]		= {inst_bytes[207][2], inst_bytes[207][3], inst_bytes[207][4], inst_bytes[207][5], inst_bytes[207][6], inst_bytes[208][0], inst_bytes[208][1], inst_bytes[208][2]};

		cache_lines[128]		= {inst_bytes[208][3], inst_bytes[208][4], inst_bytes[208][5], inst_bytes[208][6], inst_bytes[208][7], inst_bytes[209][0], inst_bytes[209][1], inst_bytes[209][2]};

		cache_lines[129]		= {inst_bytes[210][0], inst_bytes[210][1], inst_bytes[210][2], inst_bytes[211][0], inst_bytes[211][1], inst_bytes[211][2], inst_bytes[211][3], inst_bytes[212][0]};

		cache_lines[130]		= {inst_bytes[212][1], inst_bytes[212][2], inst_bytes[212][3], inst_bytes[212][4], inst_bytes[212][5], inst_bytes[212][6], inst_bytes[213][0], inst_bytes[213][1]};

		cache_lines[131]		= {inst_bytes[213][2], inst_bytes[213][3], inst_bytes[214][0], inst_bytes[214][1], inst_bytes[214][2], inst_bytes[214][3], inst_bytes[214][4], inst_bytes[215][0]};

		cache_lines[132]		= {inst_bytes[215][1], inst_bytes[215][2], inst_bytes[215][3], inst_bytes[215][4], inst_bytes[215][5], inst_bytes[215][6], inst_bytes[216][0], inst_bytes[216][1]};

		cache_lines[133]		= {inst_bytes[216][2], inst_bytes[216][3], inst_bytes[216][4], inst_bytes[216][5], inst_bytes[216][6], inst_bytes[216][7], inst_bytes[217][0], inst_bytes[217][1]};

		cache_lines[134]		= {inst_bytes[217][2], inst_bytes[218][0], inst_bytes[218][1], inst_bytes[218][2], inst_bytes[219][0], inst_bytes[219][1], inst_bytes[219][2], inst_bytes[219][3]};

		cache_lines[135]		= {inst_bytes[220][0], inst_bytes[220][1], inst_bytes[220][2], inst_bytes[220][3], inst_bytes[220][4], inst_bytes[220][5], inst_bytes[220][6], inst_bytes[221][0]};

		cache_lines[136]		= {inst_bytes[221][1], inst_bytes[221][2], inst_bytes[221][3], inst_bytes[222][0], inst_bytes[222][1], inst_bytes[222][2], inst_bytes[222][3], inst_bytes[222][4]};

		cache_lines[137]		= {inst_bytes[223][0], inst_bytes[223][1], inst_bytes[223][2], inst_bytes[223][3], inst_bytes[223][4], inst_bytes[223][5], inst_bytes[223][6], inst_bytes[224][0]};

		cache_lines[138]		= {inst_bytes[224][1], inst_bytes[224][2], inst_bytes[224][3], inst_bytes[224][4], inst_bytes[224][5], inst_bytes[224][6], inst_bytes[224][7], inst_bytes[225][0]};

		cache_lines[139]		= {inst_bytes[225][1], inst_bytes[225][2], inst_bytes[226][0], inst_bytes[226][1], inst_bytes[226][2], inst_bytes[227][0], inst_bytes[227][1], inst_bytes[227][2]};

		cache_lines[140]		= {inst_bytes[227][3], inst_bytes[228][0], inst_bytes[228][1], inst_bytes[228][2], inst_bytes[228][3], inst_bytes[228][4], inst_bytes[228][5], inst_bytes[228][6]};

		cache_lines[141]		= {inst_bytes[229][0], inst_bytes[229][1], inst_bytes[229][2], inst_bytes[229][3], inst_bytes[230][0], inst_bytes[230][1], inst_bytes[230][2], inst_bytes[230][3]};

		cache_lines[142]		= {inst_bytes[230][4], inst_bytes[231][0], inst_bytes[231][1], inst_bytes[231][2], inst_bytes[231][3], inst_bytes[231][4], inst_bytes[231][5], inst_bytes[231][6]};

		cache_lines[143]		= {inst_bytes[232][0], inst_bytes[232][1], inst_bytes[232][2], inst_bytes[232][3], inst_bytes[232][4], inst_bytes[232][5], inst_bytes[232][6], inst_bytes[232][7]};

		cache_lines[144]		= {inst_bytes[233][0], inst_bytes[233][1], inst_bytes[233][2], inst_bytes[234][0], inst_bytes[234][1], inst_bytes[234][2], inst_bytes[235][0], inst_bytes[235][1]};

		cache_lines[145]		= {inst_bytes[235][2], inst_bytes[235][3], inst_bytes[236][0], inst_bytes[236][1], inst_bytes[236][2], inst_bytes[236][3], inst_bytes[236][4], inst_bytes[236][5]};

		cache_lines[146]		= {inst_bytes[236][6], inst_bytes[237][0], inst_bytes[237][1], inst_bytes[237][2], inst_bytes[237][3], inst_bytes[238][0], inst_bytes[238][1], inst_bytes[238][2]};

		cache_lines[147]		= {inst_bytes[238][3], inst_bytes[238][4], inst_bytes[239][0], inst_bytes[239][1], inst_bytes[239][2], inst_bytes[239][3], inst_bytes[239][4], inst_bytes[239][5]};

		cache_lines[148]		= {inst_bytes[239][6], inst_bytes[240][0], inst_bytes[240][1], inst_bytes[240][2], inst_bytes[240][3], inst_bytes[240][4], inst_bytes[240][5], inst_bytes[240][6]};

		cache_lines[149]		= {inst_bytes[240][7], inst_bytes[241][0], inst_bytes[241][1], inst_bytes[241][2], inst_bytes[242][0], inst_bytes[243][0], inst_bytes[244][0], inst_bytes[244][1]};

		cache_lines[150]		= {inst_bytes[245][0], inst_bytes[245][1], inst_bytes[245][2], inst_bytes[246][0], inst_bytes[246][1], inst_bytes[246][2], inst_bytes[246][3], inst_bytes[246][4]};

		cache_lines[151]		= {inst_bytes[246][5], inst_bytes[247][0], inst_bytes[247][1], inst_bytes[247][2], inst_bytes[248][0], inst_bytes[248][1], inst_bytes[248][2], inst_bytes[248][3]};

		cache_lines[152]		= {inst_bytes[249][0], inst_bytes[249][1], inst_bytes[249][2], inst_bytes[249][3], inst_bytes[249][4], inst_bytes[249][5], inst_bytes[250][0], inst_bytes[250][1]};

		cache_lines[153]		= {inst_bytes[250][2], inst_bytes[250][3], inst_bytes[250][4], inst_bytes[250][5], inst_bytes[250][6], inst_bytes[251][0], inst_bytes[251][1], inst_bytes[252][0]};

		cache_lines[154]		= {inst_bytes[252][1], inst_bytes[253][0], inst_bytes[253][1], inst_bytes[253][2], inst_bytes[254][0], inst_bytes[254][1], inst_bytes[254][2], inst_bytes[254][3]};

		cache_lines[155]		= {inst_bytes[254][4], inst_bytes[254][5], inst_bytes[255][0], inst_bytes[255][1], inst_bytes[255][2], inst_bytes[256][0], inst_bytes[256][1], inst_bytes[256][2]};

		cache_lines[156]		= {inst_bytes[256][3], inst_bytes[257][0], inst_bytes[257][1], inst_bytes[257][2], inst_bytes[257][3], inst_bytes[257][4], inst_bytes[257][5], inst_bytes[258][0]};

		cache_lines[157]		= {inst_bytes[258][1], inst_bytes[258][2], inst_bytes[258][3], inst_bytes[258][4], inst_bytes[258][5], inst_bytes[258][6], inst_bytes[259][0], inst_bytes[259][1]};

		cache_lines[158]		= {inst_bytes[260][0], inst_bytes[260][1], inst_bytes[261][0], inst_bytes[261][1], inst_bytes[261][2], inst_bytes[262][0], inst_bytes[262][1], inst_bytes[262][2]};

		cache_lines[159]		= {inst_bytes[262][3], inst_bytes[262][4], inst_bytes[262][5], inst_bytes[263][0], inst_bytes[263][1], inst_bytes[263][2], inst_bytes[264][0], inst_bytes[264][1]};

		cache_lines[160]		= {inst_bytes[264][2], inst_bytes[264][3], inst_bytes[265][0], inst_bytes[265][1], inst_bytes[265][2], inst_bytes[265][3], inst_bytes[265][4], inst_bytes[265][5]};

		cache_lines[161]		= {inst_bytes[266][0], inst_bytes[266][1], inst_bytes[266][2], inst_bytes[266][3], inst_bytes[266][4], inst_bytes[266][5], inst_bytes[266][6], inst_bytes[267][0]};

		cache_lines[162]		= {inst_bytes[267][1], inst_bytes[268][0], inst_bytes[268][1], inst_bytes[269][0], inst_bytes[270][0], inst_bytes[271][0], inst_bytes[271][1], inst_bytes[272][0]};

		cache_lines[163]		= {inst_bytes[272][1], inst_bytes[273][0], inst_bytes[273][1], inst_bytes[273][2], inst_bytes[273][3], inst_bytes[273][4], inst_bytes[274][0], inst_bytes[274][1]};

		cache_lines[164]		= {inst_bytes[274][2], inst_bytes[274][3], inst_bytes[274][4], inst_bytes[274][5], inst_bytes[275][0], inst_bytes[275][1], inst_bytes[275][2], inst_bytes[275][3]};

		cache_lines[165]		= {inst_bytes[275][4], inst_bytes[276][0], inst_bytes[276][1], inst_bytes[276][2], inst_bytes[276][3], inst_bytes[276][4], inst_bytes[276][5], inst_bytes[277][0]};

		cache_lines[166]		= {inst_bytes[277][1], inst_bytes[278][0], inst_bytes[278][1], inst_bytes[278][2], inst_bytes[278][3], inst_bytes[279][0], inst_bytes[279][1], inst_bytes[279][2]};

		cache_lines[167]		= {inst_bytes[279][3], inst_bytes[279][4], inst_bytes[280][0], inst_bytes[280][1], inst_bytes[281][0], inst_bytes[281][1], inst_bytes[281][2], inst_bytes[282][0]};

		cache_lines[168]		= {inst_bytes[282][1], inst_bytes[282][2], inst_bytes[282][3], inst_bytes[282][4], inst_bytes[282][5], inst_bytes[283][0], inst_bytes[283][1], inst_bytes[283][2]};

		cache_lines[169]		= {inst_bytes[284][0], inst_bytes[284][1], inst_bytes[284][2], inst_bytes[284][3], inst_bytes[285][0], inst_bytes[285][1], inst_bytes[285][2], inst_bytes[285][3]};

		cache_lines[170]		= {inst_bytes[285][4], inst_bytes[285][5], inst_bytes[286][0], inst_bytes[286][1], inst_bytes[286][2], inst_bytes[286][3], inst_bytes[286][4], inst_bytes[286][5]};

		cache_lines[171]		= {inst_bytes[286][6], inst_bytes[287][0], inst_bytes[287][1], inst_bytes[288][0], inst_bytes[288][1], inst_bytes[289][0], inst_bytes[289][1], inst_bytes[289][2]};

		cache_lines[172]		= {inst_bytes[290][0], inst_bytes[290][1], inst_bytes[290][2], inst_bytes[290][3], inst_bytes[290][4], inst_bytes[290][5], inst_bytes[291][0], inst_bytes[291][1]};

		cache_lines[173]		= {inst_bytes[291][2], inst_bytes[292][0], inst_bytes[292][1], inst_bytes[292][2], inst_bytes[292][3], inst_bytes[293][0], inst_bytes[293][1], inst_bytes[293][2]};

		cache_lines[174]		= {inst_bytes[293][3], inst_bytes[293][4], inst_bytes[293][5], inst_bytes[294][0], inst_bytes[294][1], inst_bytes[294][2], inst_bytes[294][3], inst_bytes[294][4]};

		cache_lines[175]		= {inst_bytes[294][5], inst_bytes[294][6], inst_bytes[295][0], inst_bytes[295][1], inst_bytes[296][0], inst_bytes[296][1], inst_bytes[296][2], inst_bytes[296][3]};

		cache_lines[176]		= {inst_bytes[296][4], inst_bytes[296][5], inst_bytes[297][0], inst_bytes[297][1], inst_bytes[297][2], inst_bytes[297][3], inst_bytes[297][4], inst_bytes[297][5]};

		cache_lines[177]		= {inst_bytes[297][6], inst_bytes[298][0], inst_bytes[298][1], inst_bytes[299][0], inst_bytes[299][1], inst_bytes[299][2], inst_bytes[300][0], inst_bytes[300][1]};

		cache_lines[178]		= {inst_bytes[300][2], inst_bytes[300][3], inst_bytes[300][4], inst_bytes[300][5], inst_bytes[301][0], inst_bytes[301][1], inst_bytes[301][2], inst_bytes[302][0]};

		cache_lines[179]		= {inst_bytes[302][1], inst_bytes[302][2], inst_bytes[302][3], inst_bytes[303][0], inst_bytes[303][1], inst_bytes[303][2], inst_bytes[303][3], inst_bytes[303][4]};

		cache_lines[180]		= {inst_bytes[303][5], inst_bytes[304][0], inst_bytes[304][1], inst_bytes[304][2], inst_bytes[304][3], inst_bytes[304][4], inst_bytes[304][5], inst_bytes[304][6]};

		cache_lines[181]		= {inst_bytes[305][0], inst_bytes[305][1], inst_bytes[306][0], inst_bytes[306][1], inst_bytes[307][0], inst_bytes[307][1], inst_bytes[307][2], inst_bytes[308][0]};

		cache_lines[182]		= {inst_bytes[308][1], inst_bytes[308][2], inst_bytes[308][3], inst_bytes[308][4], inst_bytes[308][5], inst_bytes[309][0], inst_bytes[309][1], inst_bytes[309][2]};

		cache_lines[183]		= {inst_bytes[310][0], inst_bytes[310][1], inst_bytes[310][2], inst_bytes[310][3], inst_bytes[311][0], inst_bytes[311][1], inst_bytes[311][2], inst_bytes[311][3]};

		cache_lines[184]		= {inst_bytes[311][4], inst_bytes[311][5], inst_bytes[312][0], inst_bytes[312][1], inst_bytes[312][2], inst_bytes[312][3], inst_bytes[312][4], inst_bytes[312][5]};

		cache_lines[185]		= {inst_bytes[312][6], inst_bytes[313][0], inst_bytes[313][1], inst_bytes[314][0], inst_bytes[314][1], inst_bytes[315][0], inst_bytes[315][1], inst_bytes[315][2]};

		cache_lines[186]		= {inst_bytes[316][0], inst_bytes[316][1], inst_bytes[316][2], inst_bytes[316][3], inst_bytes[316][4], inst_bytes[316][5], inst_bytes[317][0], inst_bytes[317][1]};

		cache_lines[187]		= {inst_bytes[317][2], inst_bytes[318][0], inst_bytes[318][1], inst_bytes[318][2], inst_bytes[318][3], inst_bytes[319][0], inst_bytes[319][1], inst_bytes[319][2]};

		cache_lines[188]		= {inst_bytes[319][3], inst_bytes[319][4], inst_bytes[319][5], inst_bytes[320][0], inst_bytes[320][1], inst_bytes[320][2], inst_bytes[320][3], inst_bytes[320][4]};

		cache_lines[189]		= {inst_bytes[320][5], inst_bytes[320][6], inst_bytes[321][0], inst_bytes[321][1], inst_bytes[322][0], inst_bytes[322][1], inst_bytes[323][0], inst_bytes[323][1]};

		cache_lines[190]		= {inst_bytes[323][2], inst_bytes[324][0], inst_bytes[324][1], inst_bytes[324][2], inst_bytes[324][3], inst_bytes[324][4], inst_bytes[324][5], inst_bytes[325][0]};

		cache_lines[191]		= {inst_bytes[325][1], inst_bytes[325][2], inst_bytes[326][0], inst_bytes[326][1], inst_bytes[326][2], inst_bytes[326][3], inst_bytes[327][0], inst_bytes[327][1]};

		cache_lines[192]		= {inst_bytes[327][2], inst_bytes[327][3], inst_bytes[327][4], inst_bytes[327][5], inst_bytes[328][0], inst_bytes[328][1], inst_bytes[328][2], inst_bytes[328][3]};

		cache_lines[193]		= {inst_bytes[328][4], inst_bytes[328][5], inst_bytes[328][6], inst_bytes[329][0], inst_bytes[329][1], inst_bytes[330][0], inst_bytes[330][1], inst_bytes[331][0]};

		cache_lines[194]		= {inst_bytes[331][1], inst_bytes[331][2], inst_bytes[332][0], inst_bytes[332][1], inst_bytes[332][2], inst_bytes[332][3], inst_bytes[332][4], inst_bytes[332][5]};

		cache_lines[195]		= {inst_bytes[333][0], inst_bytes[333][1], inst_bytes[333][2], inst_bytes[334][0], inst_bytes[334][1], inst_bytes[334][2], inst_bytes[334][3], inst_bytes[335][0]};

		cache_lines[196]		= {inst_bytes[335][1], inst_bytes[335][2], inst_bytes[335][3], inst_bytes[335][4], inst_bytes[335][5], inst_bytes[336][0], inst_bytes[336][1], inst_bytes[336][2]};

		cache_lines[197]		= {inst_bytes[336][3], inst_bytes[336][4], inst_bytes[336][5], inst_bytes[336][6], inst_bytes[337][0], inst_bytes[337][1], inst_bytes[338][0], inst_bytes[338][1]};

		cache_lines[198]		= {inst_bytes[339][0], inst_bytes[339][1], inst_bytes[339][2], inst_bytes[340][0], inst_bytes[340][1], inst_bytes[340][2], inst_bytes[340][3], inst_bytes[340][4]};

		cache_lines[199]		= {inst_bytes[340][5], inst_bytes[341][0], inst_bytes[341][1], inst_bytes[341][2], inst_bytes[342][0], inst_bytes[342][1], inst_bytes[342][2], inst_bytes[342][3]};

		cache_lines[200]		= {inst_bytes[343][0], inst_bytes[343][1], inst_bytes[343][2], inst_bytes[343][3], inst_bytes[343][4], inst_bytes[343][5], inst_bytes[344][0], inst_bytes[344][1]};

		cache_lines[201]		= {inst_bytes[344][2], inst_bytes[344][3], inst_bytes[344][4], inst_bytes[344][5], inst_bytes[344][6], inst_bytes[345][0], inst_bytes[345][1], inst_bytes[346][0]};

		cache_lines[202]		= {inst_bytes[346][1], inst_bytes[347][0], inst_bytes[347][1], inst_bytes[347][2], inst_bytes[348][0], inst_bytes[348][1], inst_bytes[348][2], inst_bytes[348][3]};

		cache_lines[203]		= {inst_bytes[348][4], inst_bytes[348][5], inst_bytes[349][0], inst_bytes[349][1], inst_bytes[349][2], inst_bytes[350][0], inst_bytes[350][1], inst_bytes[350][2]};

		cache_lines[204]		= {inst_bytes[350][3], inst_bytes[351][0], inst_bytes[351][1], inst_bytes[351][2], inst_bytes[351][3], inst_bytes[351][4], inst_bytes[351][5], inst_bytes[352][0]};

		cache_lines[205]		= {inst_bytes[352][1], inst_bytes[352][2], inst_bytes[352][3], inst_bytes[352][4], inst_bytes[352][5], inst_bytes[352][6], inst_bytes[353][0], inst_bytes[353][1]};

		cache_lines[206]		= {inst_bytes[354][0], inst_bytes[354][1], inst_bytes[355][0], inst_bytes[355][1], inst_bytes[355][2], inst_bytes[356][0], inst_bytes[356][1], inst_bytes[356][2]};

		cache_lines[207]		= {inst_bytes[356][3], inst_bytes[356][4], inst_bytes[356][5], inst_bytes[357][0], inst_bytes[357][1], inst_bytes[357][2], inst_bytes[358][0], inst_bytes[358][1]};

		cache_lines[208]		= {inst_bytes[358][2], inst_bytes[358][3], inst_bytes[359][0], inst_bytes[359][1], inst_bytes[359][2], inst_bytes[359][3], inst_bytes[359][4], inst_bytes[359][5]};

		cache_lines[209]		= {inst_bytes[360][0], inst_bytes[360][1], inst_bytes[360][2], inst_bytes[360][3], inst_bytes[360][4], inst_bytes[360][5], inst_bytes[360][6], inst_bytes[361][0]};

		cache_lines[210]		= {inst_bytes[361][1], inst_bytes[362][0], inst_bytes[362][1], inst_bytes[363][0], inst_bytes[363][1], inst_bytes[363][2], inst_bytes[363][3], inst_bytes[364][0]};

		cache_lines[211]		= {inst_bytes[364][1], inst_bytes[364][2], inst_bytes[364][3], inst_bytes[364][4], inst_bytes[365][0], inst_bytes[365][1], inst_bytes[365][2], inst_bytes[366][0]};

		cache_lines[212]		= {inst_bytes[366][1], inst_bytes[366][2], inst_bytes[366][3], inst_bytes[367][0], inst_bytes[367][1], inst_bytes[367][2], inst_bytes[367][3], inst_bytes[367][4]};

		cache_lines[213]		= {inst_bytes[367][5], inst_bytes[367][6], inst_bytes[368][0], inst_bytes[368][1], inst_bytes[368][2], inst_bytes[368][3], inst_bytes[369][0], inst_bytes[369][1]};

		cache_lines[214]		= {inst_bytes[369][2], inst_bytes[369][3], inst_bytes[369][4], inst_bytes[370][0], inst_bytes[370][1], inst_bytes[370][2], inst_bytes[370][3], inst_bytes[370][4]};

		cache_lines[215]		= {inst_bytes[370][5], inst_bytes[370][6], inst_bytes[371][0], inst_bytes[371][1], inst_bytes[371][2], inst_bytes[371][3], inst_bytes[371][4], inst_bytes[371][5]};

		cache_lines[216]		= {inst_bytes[371][6], inst_bytes[371][7], inst_bytes[372][0], inst_bytes[372][1], inst_bytes[372][2], inst_bytes[373][0], inst_bytes[373][1], inst_bytes[373][2]};

		cache_lines[217]		= {inst_bytes[373][3], inst_bytes[373][4], inst_bytes[374][0], inst_bytes[374][1], inst_bytes[374][2], inst_bytes[374][3], inst_bytes[374][4], inst_bytes[374][5]};

		cache_lines[218]		= {inst_bytes[375][0], inst_bytes[375][1], inst_bytes[375][2], inst_bytes[375][3], inst_bytes[375][4], inst_bytes[375][5], inst_bytes[375][6], inst_bytes[375][7]};

		cache_lines[219]		= {inst_bytes[375][8], inst_bytes[376][0], inst_bytes[376][1], inst_bytes[376][2], inst_bytes[376][3], inst_bytes[376][4], inst_bytes[376][5], inst_bytes[377][0]};

		cache_lines[220]		= {inst_bytes[377][1], inst_bytes[377][2], inst_bytes[377][3], inst_bytes[377][4], inst_bytes[377][5], inst_bytes[377][6], inst_bytes[378][0], inst_bytes[378][1]};

		cache_lines[221]		= {inst_bytes[378][2], inst_bytes[378][3], inst_bytes[378][4], inst_bytes[378][5], inst_bytes[378][6], inst_bytes[378][7], inst_bytes[378][8], inst_bytes[379][0]};

		cache_lines[222]		= {inst_bytes[379][1], inst_bytes[379][2], inst_bytes[379][3], inst_bytes[379][4], inst_bytes[379][5], inst_bytes[379][6], inst_bytes[379][7], inst_bytes[379][8]};

		cache_lines[223]		= {inst_bytes[379][9], inst_bytes[380][0], inst_bytes[380][1], inst_bytes[380][2], inst_bytes[380][3], inst_bytes[380][4], inst_bytes[381][0], inst_bytes[381][1]};

		cache_lines[224]		= {inst_bytes[381][2], inst_bytes[381][3], inst_bytes[381][4], inst_bytes[381][5], inst_bytes[382][0], inst_bytes[382][1], inst_bytes[382][2], inst_bytes[382][3]};

		cache_lines[225]		= {inst_bytes[382][4], inst_bytes[382][5], inst_bytes[382][6], inst_bytes[383][0], inst_bytes[383][1], inst_bytes[383][2], inst_bytes[383][3], inst_bytes[383][4]};

		cache_lines[226]		= {inst_bytes[383][5], inst_bytes[383][6], inst_bytes[383][7], inst_bytes[383][8], inst_bytes[383][9], inst_bytes[384][0], inst_bytes[384][1], inst_bytes[384][2]};

		cache_lines[227]		= {inst_bytes[384][3], inst_bytes[384][4], inst_bytes[384][5], inst_bytes[384][6], inst_bytes[385][0], inst_bytes[385][1], inst_bytes[385][2], inst_bytes[385][3]};

		cache_lines[228]		= {inst_bytes[385][4], inst_bytes[385][5], inst_bytes[385][6], inst_bytes[385][7], inst_bytes[386][0], inst_bytes[386][1], inst_bytes[386][2], inst_bytes[386][3]};

		cache_lines[229]		= {inst_bytes[386][4], inst_bytes[386][5], inst_bytes[386][6], inst_bytes[386][7], inst_bytes[386][8], inst_bytes[386][9], inst_bytes[387][0], inst_bytes[387][1]};

		cache_lines[230]		= {inst_bytes[387][2], inst_bytes[387][3], inst_bytes[387][4], inst_bytes[387][5], inst_bytes[387][6], inst_bytes[387][7], inst_bytes[387][8], inst_bytes[387][9]};

		cache_lines[231]		= {inst_bytes[387][10], inst_bytes[388][0], inst_bytes[388][1], inst_bytes[388][2], inst_bytes[388][3], inst_bytes[388][4], inst_bytes[388][5], inst_bytes[389][0]};

		cache_lines[232]		= {inst_bytes[389][1], inst_bytes[389][2], inst_bytes[390][0], inst_bytes[390][1], inst_bytes[390][2], inst_bytes[390][3], inst_bytes[391][0], inst_bytes[391][1]};

		cache_lines[233]		= {inst_bytes[391][2], inst_bytes[391][3], inst_bytes[391][4], inst_bytes[391][5], inst_bytes[391][6], inst_bytes[392][0], inst_bytes[392][1], inst_bytes[392][2]};

		cache_lines[234]		= {inst_bytes[392][3], inst_bytes[393][0], inst_bytes[393][1], inst_bytes[393][2], inst_bytes[393][3], inst_bytes[393][4], inst_bytes[394][0], inst_bytes[394][1]};

		cache_lines[235]		= {inst_bytes[394][2], inst_bytes[394][3], inst_bytes[394][4], inst_bytes[394][5], inst_bytes[394][6], inst_bytes[395][0], inst_bytes[395][1], inst_bytes[395][2]};

		cache_lines[236]		= {inst_bytes[395][3], inst_bytes[395][4], inst_bytes[395][5], inst_bytes[395][6], inst_bytes[395][7], inst_bytes[396][0], inst_bytes[396][1], inst_bytes[396][2]};

		cache_lines[237]		= {inst_bytes[397][0], inst_bytes[397][1], inst_bytes[397][2], inst_bytes[398][0], inst_bytes[398][1], inst_bytes[398][2], inst_bytes[398][3], inst_bytes[399][0]};

		cache_lines[238]		= {inst_bytes[399][1], inst_bytes[399][2], inst_bytes[399][3], inst_bytes[399][4], inst_bytes[399][5], inst_bytes[399][6], inst_bytes[400][0], inst_bytes[400][1]};

		cache_lines[239]		= {inst_bytes[400][2], inst_bytes[400][3], inst_bytes[401][0], inst_bytes[401][1], inst_bytes[401][2], inst_bytes[401][3], inst_bytes[401][4], inst_bytes[402][0]};

		cache_lines[240]		= {inst_bytes[402][1], inst_bytes[402][2], inst_bytes[402][3], inst_bytes[402][4], inst_bytes[402][5], inst_bytes[402][6], inst_bytes[403][0], inst_bytes[403][1]};

		cache_lines[241]		= {inst_bytes[403][2], inst_bytes[403][3], inst_bytes[403][4], inst_bytes[403][5], inst_bytes[403][6], inst_bytes[403][7], inst_bytes[404][0], inst_bytes[404][1]};

		cache_lines[242]		= {inst_bytes[404][2], inst_bytes[405][0], inst_bytes[405][1], inst_bytes[406][0], inst_bytes[406][1], inst_bytes[406][2], inst_bytes[407][0], inst_bytes[407][1]};

		cache_lines[243]		= {inst_bytes[407][2], inst_bytes[407][3], inst_bytes[407][4], inst_bytes[407][5], inst_bytes[408][0], inst_bytes[408][1], inst_bytes[408][2], inst_bytes[409][0]};

		cache_lines[244]		= {inst_bytes[409][1], inst_bytes[409][2], inst_bytes[409][3], inst_bytes[410][0], inst_bytes[410][1], inst_bytes[410][2], inst_bytes[410][3], inst_bytes[410][4]};

		cache_lines[245]		= {inst_bytes[410][5], inst_bytes[411][0], inst_bytes[411][1], inst_bytes[411][2], inst_bytes[411][3], inst_bytes[411][4], inst_bytes[411][5], inst_bytes[411][6]};

		cache_lines[246]		= {inst_bytes[412][0], inst_bytes[412][1], inst_bytes[413][0], inst_bytes[413][1], inst_bytes[414][0], inst_bytes[414][1], inst_bytes[414][2], inst_bytes[415][0]};

		cache_lines[247]		= {inst_bytes[415][1], inst_bytes[415][2], inst_bytes[415][3], inst_bytes[415][4], inst_bytes[415][5], inst_bytes[416][0], inst_bytes[416][1], inst_bytes[416][2]};

		cache_lines[248]		= {inst_bytes[417][0], inst_bytes[417][1], inst_bytes[417][2], inst_bytes[417][3], inst_bytes[418][0], inst_bytes[418][1], inst_bytes[418][2], inst_bytes[418][3]};

		cache_lines[249]		= {inst_bytes[418][4], inst_bytes[418][5], inst_bytes[419][0], inst_bytes[419][1], inst_bytes[419][2], inst_bytes[419][3], inst_bytes[419][4], inst_bytes[419][5]};

		cache_lines[250]		= {inst_bytes[419][6], inst_bytes[420][0], inst_bytes[420][1], inst_bytes[421][0], inst_bytes[421][1], inst_bytes[422][0], inst_bytes[422][1], inst_bytes[422][2]};

		cache_lines[251]		= {inst_bytes[423][0], inst_bytes[423][1], inst_bytes[423][2], inst_bytes[423][3], inst_bytes[423][4], inst_bytes[423][5], inst_bytes[424][0], inst_bytes[424][1]};

		cache_lines[252]		= {inst_bytes[424][2], inst_bytes[425][0], inst_bytes[425][1], inst_bytes[425][2], inst_bytes[425][3], inst_bytes[426][0], inst_bytes[426][1], inst_bytes[426][2]};

		cache_lines[253]		= {inst_bytes[426][3], inst_bytes[426][4], inst_bytes[426][5], inst_bytes[427][0], inst_bytes[427][1], inst_bytes[427][2], inst_bytes[427][3], inst_bytes[427][4]};

		cache_lines[254]		= {inst_bytes[427][5], inst_bytes[427][6], inst_bytes[428][0], inst_bytes[428][1], inst_bytes[429][0], inst_bytes[429][1], inst_bytes[430][0], inst_bytes[430][1]};

		cache_lines[255]		= {inst_bytes[430][2], inst_bytes[430][3], inst_bytes[431][0], inst_bytes[431][1], inst_bytes[431][2], inst_bytes[431][3], inst_bytes[431][4], inst_bytes[432][0]};

		cache_lines[256]		= {inst_bytes[432][1], inst_bytes[432][2], inst_bytes[433][0], inst_bytes[433][1], inst_bytes[433][2], inst_bytes[433][3], inst_bytes[434][0], inst_bytes[434][1]};

		cache_lines[257]		= {inst_bytes[434][2], inst_bytes[434][3], inst_bytes[434][4], inst_bytes[434][5], inst_bytes[434][6], inst_bytes[435][0], inst_bytes[435][1], inst_bytes[435][2]};

		cache_lines[258]		= {inst_bytes[435][3], inst_bytes[436][0], inst_bytes[436][1], inst_bytes[436][2], inst_bytes[436][3], inst_bytes[436][4], inst_bytes[437][0], inst_bytes[437][1]};

		cache_lines[259]		= {inst_bytes[437][2], inst_bytes[437][3], inst_bytes[437][4], inst_bytes[437][5], inst_bytes[437][6], inst_bytes[438][0], inst_bytes[438][1], inst_bytes[438][2]};

		cache_lines[260]		= {inst_bytes[438][3], inst_bytes[438][4], inst_bytes[438][5], inst_bytes[438][6], inst_bytes[438][7], inst_bytes[439][0], inst_bytes[439][1], inst_bytes[439][2]};

		cache_lines[261]		= {inst_bytes[440][0], inst_bytes[440][1], inst_bytes[440][2], inst_bytes[440][3], inst_bytes[440][4], inst_bytes[441][0], inst_bytes[441][1], inst_bytes[441][2]};

		cache_lines[262]		= {inst_bytes[441][3], inst_bytes[441][4], inst_bytes[441][5], inst_bytes[442][0], inst_bytes[442][1], inst_bytes[442][2], inst_bytes[442][3], inst_bytes[442][4]};

		cache_lines[263]		= {inst_bytes[442][5], inst_bytes[442][6], inst_bytes[442][7], inst_bytes[442][8], inst_bytes[443][0], inst_bytes[443][1], inst_bytes[443][2], inst_bytes[443][3]};

		cache_lines[264]		= {inst_bytes[443][4], inst_bytes[443][5], inst_bytes[444][0], inst_bytes[444][1], inst_bytes[444][2], inst_bytes[444][3], inst_bytes[444][4], inst_bytes[444][5]};

		cache_lines[265]		= {inst_bytes[444][6], inst_bytes[445][0], inst_bytes[445][1], inst_bytes[445][2], inst_bytes[445][3], inst_bytes[445][4], inst_bytes[445][5], inst_bytes[445][6]};

		cache_lines[266]		= {inst_bytes[445][7], inst_bytes[445][8], inst_bytes[446][0], inst_bytes[446][1], inst_bytes[446][2], inst_bytes[446][3], inst_bytes[446][4], inst_bytes[446][5]};

		cache_lines[267]		= {inst_bytes[446][6], inst_bytes[446][7], inst_bytes[446][8], inst_bytes[446][9], inst_bytes[447][0], inst_bytes[447][1], inst_bytes[447][2], inst_bytes[447][3]};

		cache_lines[268]		= {inst_bytes[447][4], inst_bytes[448][0], inst_bytes[448][1], inst_bytes[448][2], inst_bytes[448][3], inst_bytes[448][4], inst_bytes[448][5], inst_bytes[449][0]};

		cache_lines[269]		= {inst_bytes[449][1], inst_bytes[449][2], inst_bytes[449][3], inst_bytes[449][4], inst_bytes[449][5], inst_bytes[449][6], inst_bytes[450][0], inst_bytes[450][1]};

		cache_lines[270]		= {inst_bytes[450][2], inst_bytes[450][3], inst_bytes[450][4], inst_bytes[450][5], inst_bytes[450][6], inst_bytes[450][7], inst_bytes[450][8], inst_bytes[450][9]};

		cache_lines[271]		= {inst_bytes[451][0], inst_bytes[451][1], inst_bytes[451][2], inst_bytes[451][3], inst_bytes[451][4], inst_bytes[451][5], inst_bytes[451][6], inst_bytes[452][0]};

		cache_lines[272]		= {inst_bytes[452][1], inst_bytes[452][2], inst_bytes[452][3], inst_bytes[452][4], inst_bytes[452][5], inst_bytes[452][6], inst_bytes[452][7], inst_bytes[453][0]};

		cache_lines[273]		= {inst_bytes[453][1], inst_bytes[453][2], inst_bytes[453][3], inst_bytes[453][4], inst_bytes[453][5], inst_bytes[453][6], inst_bytes[453][7], inst_bytes[453][8]};

		cache_lines[274]		= {inst_bytes[453][9], inst_bytes[454][0], inst_bytes[454][1], inst_bytes[454][2], inst_bytes[454][3], inst_bytes[454][4], inst_bytes[454][5], inst_bytes[454][6]};

		cache_lines[275]		= {inst_bytes[454][7], inst_bytes[454][8], inst_bytes[454][9], inst_bytes[454][10], inst_bytes[455][0], inst_bytes[455][1], inst_bytes[455][2], inst_bytes[455][3]};

		cache_lines[276]		= {inst_bytes[455][4], inst_bytes[455][5], inst_bytes[456][0], inst_bytes[456][1], inst_bytes[456][2], inst_bytes[457][0], inst_bytes[457][1], inst_bytes[457][2]};

		cache_lines[277]		= {inst_bytes[457][3], inst_bytes[458][0], inst_bytes[458][1], inst_bytes[458][2], inst_bytes[458][3], inst_bytes[458][4], inst_bytes[458][5], inst_bytes[458][6]};

		cache_lines[278]		= {inst_bytes[459][0], inst_bytes[459][1], inst_bytes[459][2], inst_bytes[459][3], inst_bytes[460][0], inst_bytes[460][1], inst_bytes[460][2], inst_bytes[460][3]};

		cache_lines[279]		= {inst_bytes[460][4], inst_bytes[461][0], inst_bytes[461][1], inst_bytes[461][2], inst_bytes[461][3], inst_bytes[461][4], inst_bytes[461][5], inst_bytes[461][6]};

		cache_lines[280]		= {inst_bytes[462][0], inst_bytes[462][1], inst_bytes[462][2], inst_bytes[462][3], inst_bytes[462][4], inst_bytes[462][5], inst_bytes[462][6], inst_bytes[462][7]};

		cache_lines[281]		= {inst_bytes[463][0], inst_bytes[463][1], inst_bytes[463][2], inst_bytes[464][0], inst_bytes[464][1], inst_bytes[464][2], inst_bytes[465][0], inst_bytes[465][1]};

		cache_lines[282]		= {inst_bytes[465][2], inst_bytes[465][3], inst_bytes[466][0], inst_bytes[466][1], inst_bytes[466][2], inst_bytes[466][3], inst_bytes[466][4], inst_bytes[466][5]};

		cache_lines[283]		= {inst_bytes[466][6], inst_bytes[467][0], inst_bytes[467][1], inst_bytes[467][2], inst_bytes[467][3], inst_bytes[468][0], inst_bytes[468][1], inst_bytes[468][2]};

		cache_lines[284]		= {inst_bytes[468][3], inst_bytes[468][4], inst_bytes[469][0], inst_bytes[469][1], inst_bytes[469][2], inst_bytes[469][3], inst_bytes[469][4], inst_bytes[469][5]};

		cache_lines[285]		= {inst_bytes[469][6], inst_bytes[470][0], inst_bytes[470][1], inst_bytes[470][2], inst_bytes[470][3], inst_bytes[470][4], inst_bytes[470][5], inst_bytes[470][6]};

		cache_lines[286]		= {inst_bytes[470][7], inst_bytes[471][0], inst_bytes[471][1], inst_bytes[471][2], inst_bytes[472][0], inst_bytes[472][1], inst_bytes[473][0], inst_bytes[473][1]};

		cache_lines[287]		= {inst_bytes[473][2], inst_bytes[474][0], inst_bytes[474][1], inst_bytes[474][2], inst_bytes[474][3], inst_bytes[474][4], inst_bytes[474][5], inst_bytes[475][0]};

		cache_lines[288]		= {inst_bytes[475][1], inst_bytes[475][2], inst_bytes[476][0], inst_bytes[476][1], inst_bytes[476][2], inst_bytes[476][3], inst_bytes[477][0], inst_bytes[477][1]};

		cache_lines[289]		= {inst_bytes[477][2], inst_bytes[477][3], inst_bytes[477][4], inst_bytes[477][5], inst_bytes[478][0], inst_bytes[478][1], inst_bytes[478][2], inst_bytes[478][3]};

		cache_lines[290]		= {inst_bytes[478][4], inst_bytes[478][5], inst_bytes[478][6], inst_bytes[479][0], inst_bytes[479][1], inst_bytes[480][0], inst_bytes[480][1], inst_bytes[481][0]};

		cache_lines[291]		= {inst_bytes[481][1], inst_bytes[481][2], inst_bytes[482][0], inst_bytes[482][1], inst_bytes[482][2], inst_bytes[482][3], inst_bytes[482][4], inst_bytes[482][5]};

		cache_lines[292]		= {inst_bytes[483][0], inst_bytes[483][1], inst_bytes[483][2], inst_bytes[484][0], inst_bytes[484][1], inst_bytes[484][2], inst_bytes[484][3], inst_bytes[485][0]};

		cache_lines[293]		= {inst_bytes[485][1], inst_bytes[485][2], inst_bytes[485][3], inst_bytes[485][4], inst_bytes[485][5], inst_bytes[486][0], inst_bytes[486][1], inst_bytes[486][2]};

		cache_lines[294]		= {inst_bytes[486][3], inst_bytes[486][4], inst_bytes[486][5], inst_bytes[486][6], inst_bytes[487][0], inst_bytes[487][1], inst_bytes[488][0], inst_bytes[488][1]};

		cache_lines[295]		= {inst_bytes[489][0], inst_bytes[489][1], inst_bytes[489][2], inst_bytes[490][0], inst_bytes[490][1], inst_bytes[490][2], inst_bytes[490][3], inst_bytes[490][4]};

		cache_lines[296]		= {inst_bytes[490][5], inst_bytes[491][0], inst_bytes[491][1], inst_bytes[491][2], inst_bytes[492][0], inst_bytes[492][1], inst_bytes[492][2], inst_bytes[492][3]};

		cache_lines[297]		= {inst_bytes[493][0], inst_bytes[493][1], inst_bytes[493][2], inst_bytes[493][3], inst_bytes[493][4], inst_bytes[493][5], inst_bytes[494][0], inst_bytes[494][1]};

		cache_lines[298]		= {inst_bytes[494][2], inst_bytes[494][3], inst_bytes[494][4], inst_bytes[494][5], inst_bytes[494][6], inst_bytes[495][0], inst_bytes[495][1], inst_bytes[496][0]};

		cache_lines[299]		= {inst_bytes[496][1], inst_bytes[497][0], inst_bytes[497][1], inst_bytes[497][2], inst_bytes[498][0], inst_bytes[498][1], inst_bytes[498][2], inst_bytes[498][3]};

		cache_lines[300]		= {inst_bytes[498][4], inst_bytes[498][5], inst_bytes[499][0], inst_bytes[499][1], inst_bytes[499][2], inst_bytes[500][0], inst_bytes[500][1], inst_bytes[500][2]};

		cache_lines[301]		= {inst_bytes[500][3], inst_bytes[501][0], inst_bytes[501][1], inst_bytes[501][2], inst_bytes[501][3], inst_bytes[501][4], inst_bytes[501][5], inst_bytes[502][0]};

		cache_lines[302]		= {inst_bytes[502][1], inst_bytes[502][2], inst_bytes[502][3], inst_bytes[502][4], inst_bytes[502][5], inst_bytes[502][6], inst_bytes[503][0], inst_bytes[503][1]};

		cache_lines[303]		= {inst_bytes[504][0], inst_bytes[504][1], inst_bytes[505][0], inst_bytes[505][1], inst_bytes[505][2], inst_bytes[506][0], inst_bytes[506][1], inst_bytes[506][2]};

		cache_lines[304]		= {inst_bytes[506][3], inst_bytes[506][4], inst_bytes[506][5], inst_bytes[507][0], inst_bytes[507][1], inst_bytes[507][2], inst_bytes[508][0], inst_bytes[508][1]};

		cache_lines[305]		= {inst_bytes[508][2], inst_bytes[508][3], inst_bytes[509][0], inst_bytes[509][1], inst_bytes[509][2], inst_bytes[509][3], inst_bytes[509][4], inst_bytes[509][5]};

		cache_lines[306]		= {inst_bytes[510][0], inst_bytes[510][1], inst_bytes[510][2], inst_bytes[510][3], inst_bytes[510][4], inst_bytes[510][5], inst_bytes[510][6], inst_bytes[511][0]};

		cache_lines[307]		= {inst_bytes[511][1], inst_bytes[512][0], inst_bytes[512][1], inst_bytes[513][0], inst_bytes[513][1], inst_bytes[513][2], inst_bytes[514][0], inst_bytes[514][1]};

		cache_lines[308]		= {inst_bytes[514][2], inst_bytes[514][3], inst_bytes[514][4], inst_bytes[514][5], inst_bytes[515][0], inst_bytes[515][1], inst_bytes[515][2], inst_bytes[516][0]};

		cache_lines[309]		= {inst_bytes[516][1], inst_bytes[516][2], inst_bytes[516][3], inst_bytes[517][0], inst_bytes[517][1], inst_bytes[517][2], inst_bytes[517][3], inst_bytes[517][4]};

		cache_lines[310]		= {inst_bytes[517][5], inst_bytes[518][0], inst_bytes[518][1], inst_bytes[518][2], inst_bytes[518][3], inst_bytes[518][4], inst_bytes[518][5], inst_bytes[518][6]};

		cache_lines[311]		= {inst_bytes[519][0], inst_bytes[519][1], inst_bytes[520][0], inst_bytes[520][1], inst_bytes[520][2], inst_bytes[521][0], inst_bytes[521][1], inst_bytes[521][2]};

		cache_lines[312]		= {inst_bytes[521][3], inst_bytes[522][0], inst_bytes[522][1], inst_bytes[522][2], inst_bytes[522][3], inst_bytes[522][4], inst_bytes[522][5], inst_bytes[522][6]};

		cache_lines[313]		= {inst_bytes[523][0], inst_bytes[523][1], inst_bytes[523][2], inst_bytes[523][3], inst_bytes[524][0], inst_bytes[524][1], inst_bytes[524][2], inst_bytes[524][3]};

		cache_lines[314]		= {inst_bytes[524][4], inst_bytes[525][0], inst_bytes[525][1], inst_bytes[525][2], inst_bytes[525][3], inst_bytes[525][4], inst_bytes[525][5], inst_bytes[525][6]};

		cache_lines[315]		= {inst_bytes[526][0], inst_bytes[526][1], inst_bytes[526][2], inst_bytes[526][3], inst_bytes[526][4], inst_bytes[526][5], inst_bytes[526][6], inst_bytes[526][7]};

		cache_lines[316]		= {inst_bytes[527][0], inst_bytes[527][1], inst_bytes[527][2], inst_bytes[528][0], inst_bytes[528][1], inst_bytes[528][2], inst_bytes[529][0], inst_bytes[529][1]};

		cache_lines[317]		= {inst_bytes[529][2], inst_bytes[529][3], inst_bytes[530][0], inst_bytes[530][1], inst_bytes[530][2], inst_bytes[530][3], inst_bytes[530][4], inst_bytes[530][5]};

		cache_lines[318]		= {inst_bytes[530][6], inst_bytes[531][0], inst_bytes[531][1], inst_bytes[531][2], inst_bytes[531][3], inst_bytes[532][0], inst_bytes[532][1], inst_bytes[532][2]};

		cache_lines[319]		= {inst_bytes[532][3], inst_bytes[532][4], inst_bytes[533][0], inst_bytes[533][1], inst_bytes[533][2], inst_bytes[533][3], inst_bytes[533][4], inst_bytes[533][5]};

		cache_lines[320]		= {inst_bytes[533][6], inst_bytes[534][0], inst_bytes[534][1], inst_bytes[534][2], inst_bytes[534][3], inst_bytes[534][4], inst_bytes[534][5], inst_bytes[534][6]};

		cache_lines[321]		= {inst_bytes[534][7], inst_bytes[535][0], inst_bytes[535][1], inst_bytes[535][2], inst_bytes[536][0], inst_bytes[536][1], inst_bytes[536][2], inst_bytes[537][0]};

		cache_lines[322]		= {inst_bytes[537][1], inst_bytes[537][2], inst_bytes[537][3], inst_bytes[538][0], inst_bytes[538][1], inst_bytes[538][2], inst_bytes[538][3], inst_bytes[538][4]};

		cache_lines[323]		= {inst_bytes[538][5], inst_bytes[538][6], inst_bytes[539][0], inst_bytes[539][1], inst_bytes[539][2], inst_bytes[539][3], inst_bytes[540][0], inst_bytes[540][1]};

		cache_lines[324]		= {inst_bytes[540][2], inst_bytes[540][3], inst_bytes[540][4], inst_bytes[541][0], inst_bytes[541][1], inst_bytes[541][2], inst_bytes[541][3], inst_bytes[541][4]};

		cache_lines[325]		= {inst_bytes[541][5], inst_bytes[541][6], inst_bytes[542][0], inst_bytes[542][1], inst_bytes[542][2], inst_bytes[542][3], inst_bytes[542][4], inst_bytes[542][5]};

		cache_lines[326]		= {inst_bytes[542][6], inst_bytes[542][7], inst_bytes[543][0], inst_bytes[543][1], inst_bytes[543][2], inst_bytes[544][0], inst_bytes[544][1], inst_bytes[545][0]};

		cache_lines[327]		= {inst_bytes[545][1], inst_bytes[545][2], inst_bytes[546][0], inst_bytes[546][1], inst_bytes[546][2], inst_bytes[546][3], inst_bytes[546][4], inst_bytes[546][5]};

		cache_lines[328]		= {inst_bytes[547][0], inst_bytes[547][1], inst_bytes[547][2], inst_bytes[548][0], inst_bytes[548][1], inst_bytes[548][2], inst_bytes[548][3], inst_bytes[549][0]};

		cache_lines[329]		= {inst_bytes[549][1], inst_bytes[549][2], inst_bytes[549][3], inst_bytes[549][4], inst_bytes[549][5], inst_bytes[550][0], inst_bytes[550][1], inst_bytes[550][2]};

		cache_lines[330]		= {inst_bytes[550][3], inst_bytes[550][4], inst_bytes[550][5], inst_bytes[550][6], inst_bytes[551][0], inst_bytes[551][1], inst_bytes[552][0], inst_bytes[552][1]};

		cache_lines[331]		= {inst_bytes[553][0], inst_bytes[553][1], inst_bytes[553][2], inst_bytes[554][0], inst_bytes[554][1], inst_bytes[554][2], inst_bytes[554][3], inst_bytes[554][4]};

		cache_lines[332]		= {inst_bytes[554][5], inst_bytes[555][0], inst_bytes[555][1], inst_bytes[555][2], inst_bytes[556][0], inst_bytes[556][1], inst_bytes[556][2], inst_bytes[556][3]};

		cache_lines[333]		= {inst_bytes[557][0], inst_bytes[557][1], inst_bytes[557][2], inst_bytes[557][3], inst_bytes[557][4], inst_bytes[557][5], inst_bytes[558][0], inst_bytes[558][1]};

		cache_lines[334]		= {inst_bytes[558][2], inst_bytes[558][3], inst_bytes[558][4], inst_bytes[558][5], inst_bytes[558][6], inst_bytes[559][0], inst_bytes[559][1], inst_bytes[560][0]};

		cache_lines[335]		= {inst_bytes[560][1], inst_bytes[561][0], inst_bytes[562][0], inst_bytes[563][0], inst_bytes[564][0], inst_bytes[565][0], inst_bytes[565][1], inst_bytes[566][0]};

		cache_lines[336]		= {inst_bytes[566][1], inst_bytes[567][0], inst_bytes[567][1], inst_bytes[567][2], inst_bytes[567][3], inst_bytes[568][0], inst_bytes[568][1], inst_bytes[568][2]};

		cache_lines[337]		= {inst_bytes[568][3], inst_bytes[568][4], inst_bytes[569][0], inst_bytes[569][1], inst_bytes[569][2], inst_bytes[569][3], inst_bytes[569][4], inst_bytes[569][5]};

		cache_lines[338]		= {inst_bytes[569][6], inst_bytes[569][7], inst_bytes[570][0], inst_bytes[570][1], inst_bytes[570][2], inst_bytes[570][3], inst_bytes[570][4], inst_bytes[571][0]};

		cache_lines[339]		= {inst_bytes[571][1], inst_bytes[571][2], inst_bytes[571][3], inst_bytes[571][4], inst_bytes[571][5], inst_bytes[572][0], inst_bytes[572][1], inst_bytes[572][2]};

		cache_lines[340]		= {inst_bytes[572][3], inst_bytes[572][4], inst_bytes[572][5], inst_bytes[572][6], inst_bytes[572][7], inst_bytes[573][0], inst_bytes[573][1], inst_bytes[573][2]};

		cache_lines[341]		= {inst_bytes[573][3], inst_bytes[573][4], inst_bytes[573][5], inst_bytes[573][6], inst_bytes[573][7], inst_bytes[573][8], inst_bytes[574][0], inst_bytes[574][1]};

		cache_lines[342]		= {inst_bytes[574][2], inst_bytes[574][3], inst_bytes[575][0], inst_bytes[575][1], inst_bytes[576][0], inst_bytes[576][1], inst_bytes[576][2], inst_bytes[577][0]};

		cache_lines[343]		= {inst_bytes[577][1], inst_bytes[577][2], inst_bytes[577][3], inst_bytes[577][4], inst_bytes[577][5], inst_bytes[578][0], inst_bytes[578][1], inst_bytes[578][2]};

		cache_lines[344]		= {inst_bytes[579][0], inst_bytes[579][1], inst_bytes[579][2], inst_bytes[579][3], inst_bytes[580][0], inst_bytes[580][1], inst_bytes[580][2], inst_bytes[580][3]};

		cache_lines[345]		= {inst_bytes[580][4], inst_bytes[580][5], inst_bytes[581][0], inst_bytes[581][1], inst_bytes[581][2], inst_bytes[581][3], inst_bytes[581][4], inst_bytes[581][5]};

		cache_lines[346]		= {inst_bytes[581][6], inst_bytes[582][0], inst_bytes[582][1], inst_bytes[583][0], inst_bytes[583][1], inst_bytes[584][0], inst_bytes[584][1], inst_bytes[584][2]};

		cache_lines[347]		= {inst_bytes[585][0], inst_bytes[585][1], inst_bytes[585][2], inst_bytes[585][3], inst_bytes[585][4], inst_bytes[585][5], inst_bytes[586][0], inst_bytes[586][1]};

		cache_lines[348]		= {inst_bytes[586][2], inst_bytes[587][0], inst_bytes[587][1], inst_bytes[587][2], inst_bytes[587][3], inst_bytes[588][0], inst_bytes[588][1], inst_bytes[588][2]};

		cache_lines[349]		= {inst_bytes[588][3], inst_bytes[588][4], inst_bytes[588][5], inst_bytes[589][0], inst_bytes[589][1], inst_bytes[589][2], inst_bytes[589][3], inst_bytes[589][4]};

		cache_lines[350]		= {inst_bytes[589][5], inst_bytes[589][6], inst_bytes[590][0], inst_bytes[590][1], inst_bytes[591][0], inst_bytes[591][1], inst_bytes[592][0], inst_bytes[593][0]};

		cache_lines[351]		= {inst_bytes[593][1], inst_bytes[594][0], inst_bytes[594][1], inst_bytes[594][2], inst_bytes[594][3], inst_bytes[595][0], inst_bytes[595][1], inst_bytes[595][2]};

		cache_lines[352]		= {inst_bytes[595][3], inst_bytes[595][4], inst_bytes[596][0], inst_bytes[597][0], inst_bytes[598][0], inst_bytes[599][0], inst_bytes[600][0], inst_bytes[600][1]};

		cache_lines[353]		= {inst_bytes[601][0], inst_bytes[601][1], inst_bytes[602][0], inst_bytes[603][0], inst_bytes[604][0], inst_bytes[605][0], inst_bytes[606][0], inst_bytes[607][0]};

		cache_lines[354]		= {inst_bytes[607][1], inst_bytes[607][2], inst_bytes[607][3], inst_bytes[608][0], inst_bytes[608][1], inst_bytes[608][2], inst_bytes[608][3], inst_bytes[609][0]};

		cache_lines[355]		= {inst_bytes[609][1], inst_bytes[610][0], inst_bytes[610][1], inst_bytes[610][2], inst_bytes[611][0], inst_bytes[611][1], inst_bytes[611][2], inst_bytes[611][3]};

		cache_lines[356]		= {inst_bytes[611][4], inst_bytes[611][5], inst_bytes[612][0], inst_bytes[612][1], inst_bytes[612][2], inst_bytes[613][0], inst_bytes[613][1], inst_bytes[613][2]};

		cache_lines[357]		= {inst_bytes[613][3], inst_bytes[614][0], inst_bytes[614][1], inst_bytes[614][2], inst_bytes[614][3], inst_bytes[614][4], inst_bytes[614][5], inst_bytes[615][0]};

		cache_lines[358]		= {inst_bytes[615][1], inst_bytes[615][2], inst_bytes[615][3], inst_bytes[615][4], inst_bytes[615][5], inst_bytes[615][6], inst_bytes[616][0], inst_bytes[616][1]};

		cache_lines[359]		= {inst_bytes[617][0], inst_bytes[617][1], inst_bytes[618][0], inst_bytes[618][1], inst_bytes[618][2], inst_bytes[619][0], inst_bytes[619][1], inst_bytes[619][2]};

		cache_lines[360]		= {inst_bytes[619][3], inst_bytes[619][4], inst_bytes[619][5], inst_bytes[620][0], inst_bytes[620][1], inst_bytes[620][2], inst_bytes[621][0], inst_bytes[621][1]};

		cache_lines[361]		= {inst_bytes[621][2], inst_bytes[621][3], inst_bytes[622][0], inst_bytes[622][1], inst_bytes[622][2], inst_bytes[622][3], inst_bytes[622][4], inst_bytes[622][5]};

		cache_lines[362]		= {inst_bytes[623][0], inst_bytes[623][1], inst_bytes[623][2], inst_bytes[623][3], inst_bytes[623][4], inst_bytes[623][5], inst_bytes[623][6], inst_bytes[624][0]};

		cache_lines[363]		= {inst_bytes[624][1], inst_bytes[625][0], inst_bytes[625][1], inst_bytes[625][2], inst_bytes[626][0], inst_bytes[626][1], inst_bytes[626][2], inst_bytes[626][3]};

		cache_lines[364]		= {inst_bytes[627][0], inst_bytes[627][1], inst_bytes[627][2], inst_bytes[627][3], inst_bytes[627][4], inst_bytes[627][5], inst_bytes[627][6], inst_bytes[628][0]};

		cache_lines[365]		= {inst_bytes[628][1], inst_bytes[628][2], inst_bytes[628][3], inst_bytes[629][0], inst_bytes[629][1], inst_bytes[629][2], inst_bytes[629][3], inst_bytes[629][4]};

		cache_lines[366]		= {inst_bytes[630][0], inst_bytes[630][1], inst_bytes[630][2], inst_bytes[630][3], inst_bytes[630][4], inst_bytes[630][5], inst_bytes[630][6], inst_bytes[631][0]};

		cache_lines[367]		= {inst_bytes[631][1], inst_bytes[631][2], inst_bytes[631][3], inst_bytes[631][4], inst_bytes[631][5], inst_bytes[631][6], inst_bytes[631][7], inst_bytes[632][0]};

		cache_lines[368]		= {inst_bytes[632][1], inst_bytes[632][2], inst_bytes[633][0], inst_bytes[633][1], inst_bytes[634][0], inst_bytes[634][1], inst_bytes[634][2], inst_bytes[635][0]};

		cache_lines[369]		= {inst_bytes[635][1], inst_bytes[635][2], inst_bytes[635][3], inst_bytes[635][4], inst_bytes[635][5], inst_bytes[636][0], inst_bytes[636][1], inst_bytes[636][2]};

		cache_lines[370]		= {inst_bytes[637][0], inst_bytes[637][1], inst_bytes[637][2], inst_bytes[637][3], inst_bytes[638][0], inst_bytes[638][1], inst_bytes[638][2], inst_bytes[638][3]};

		cache_lines[371]		= {inst_bytes[638][4], inst_bytes[638][5], inst_bytes[639][0], inst_bytes[639][1], inst_bytes[639][2], inst_bytes[639][3], inst_bytes[639][4], inst_bytes[639][5]};

		cache_lines[372]		= {inst_bytes[639][6], inst_bytes[640][0], inst_bytes[640][1], inst_bytes[641][0], inst_bytes[641][1], inst_bytes[642][0], inst_bytes[642][1], inst_bytes[642][2]};

		cache_lines[373]		= {inst_bytes[643][0], inst_bytes[643][1], inst_bytes[643][2], inst_bytes[643][3], inst_bytes[643][4], inst_bytes[643][5], inst_bytes[644][0], inst_bytes[644][1]};

		cache_lines[374]		= {inst_bytes[644][2], inst_bytes[645][0], inst_bytes[645][1], inst_bytes[645][2], inst_bytes[645][3], inst_bytes[646][0], inst_bytes[646][1], inst_bytes[646][2]};

		cache_lines[375]		= {inst_bytes[646][3], inst_bytes[646][4], inst_bytes[646][5], inst_bytes[647][0], inst_bytes[647][1], inst_bytes[647][2], inst_bytes[647][3], inst_bytes[647][4]};

		cache_lines[376]		= {inst_bytes[647][5], inst_bytes[647][6], inst_bytes[648][0], inst_bytes[648][1], inst_bytes[649][0], inst_bytes[649][1], inst_bytes[649][2], inst_bytes[650][0]};

		cache_lines[377]		= {inst_bytes[650][1], inst_bytes[650][2], inst_bytes[650][3], inst_bytes[651][0], inst_bytes[651][1], inst_bytes[651][2], inst_bytes[651][3], inst_bytes[651][4]};

		cache_lines[378]		= {inst_bytes[651][5], inst_bytes[651][6], inst_bytes[652][0], inst_bytes[652][1], inst_bytes[652][2], inst_bytes[652][3], inst_bytes[653][0], inst_bytes[653][1]};

		cache_lines[379]		= {inst_bytes[653][2], inst_bytes[653][3], inst_bytes[653][4], inst_bytes[654][0], inst_bytes[654][1], inst_bytes[654][2], inst_bytes[654][3], inst_bytes[654][4]};

		cache_lines[380]		= {inst_bytes[654][5], inst_bytes[654][6], inst_bytes[655][0], inst_bytes[655][1], inst_bytes[655][2], inst_bytes[655][3], inst_bytes[655][4], inst_bytes[655][5]};

		cache_lines[381]		= {inst_bytes[655][6], inst_bytes[655][7], inst_bytes[656][0], inst_bytes[656][1], inst_bytes[656][2], inst_bytes[657][0], inst_bytes[657][1], inst_bytes[658][0]};

		cache_lines[382]		= {inst_bytes[658][1], inst_bytes[658][2], inst_bytes[659][0], inst_bytes[659][1], inst_bytes[659][2], inst_bytes[659][3], inst_bytes[659][4], inst_bytes[659][5]};

		cache_lines[383]		= {inst_bytes[660][0], inst_bytes[660][1], inst_bytes[660][2], inst_bytes[661][0], inst_bytes[661][1], inst_bytes[661][2], inst_bytes[661][3], inst_bytes[662][0]};

		cache_lines[384]		= {inst_bytes[662][1], inst_bytes[662][2], inst_bytes[662][3], inst_bytes[662][4], inst_bytes[662][5], inst_bytes[663][0], inst_bytes[663][1], inst_bytes[663][2]};

		cache_lines[385]		= {inst_bytes[663][3], inst_bytes[663][4], inst_bytes[663][5], inst_bytes[663][6], inst_bytes[664][0], inst_bytes[664][1], inst_bytes[665][0], inst_bytes[665][1]};

		cache_lines[386]		= {inst_bytes[666][0], inst_bytes[666][1], inst_bytes[666][2], inst_bytes[667][0], inst_bytes[667][1], inst_bytes[667][2], inst_bytes[667][3], inst_bytes[667][4]};

		cache_lines[387]		= {inst_bytes[667][5], inst_bytes[668][0], inst_bytes[668][1], inst_bytes[668][2], inst_bytes[669][0], inst_bytes[669][1], inst_bytes[669][2], inst_bytes[669][3]};

		cache_lines[388]		= {inst_bytes[670][0], inst_bytes[670][1], inst_bytes[670][2], inst_bytes[670][3], inst_bytes[670][4], inst_bytes[670][5], inst_bytes[671][0], inst_bytes[671][1]};

		cache_lines[389]		= {inst_bytes[671][2], inst_bytes[671][3], inst_bytes[671][4], inst_bytes[671][5], inst_bytes[671][6], inst_bytes[672][0], inst_bytes[672][1], inst_bytes[673][0]};

		cache_lines[390]		= {inst_bytes[673][1], inst_bytes[673][2], inst_bytes[674][0], inst_bytes[674][1], inst_bytes[674][2], inst_bytes[674][3], inst_bytes[675][0], inst_bytes[675][1]};

		cache_lines[391]		= {inst_bytes[675][2], inst_bytes[675][3], inst_bytes[675][4], inst_bytes[675][5], inst_bytes[675][6], inst_bytes[676][0], inst_bytes[676][1], inst_bytes[676][2]};

		cache_lines[392]		= {inst_bytes[676][3], inst_bytes[677][0], inst_bytes[677][1], inst_bytes[677][2], inst_bytes[677][3], inst_bytes[677][4], inst_bytes[678][0], inst_bytes[678][1]};

		cache_lines[393]		= {inst_bytes[678][2], inst_bytes[678][3], inst_bytes[678][4], inst_bytes[678][5], inst_bytes[678][6], inst_bytes[679][0], inst_bytes[679][1], inst_bytes[679][2]};

		cache_lines[394]		= {inst_bytes[679][3], inst_bytes[679][4], inst_bytes[679][5], inst_bytes[679][6], inst_bytes[679][7], inst_bytes[680][0], inst_bytes[680][1], inst_bytes[680][2]};

		cache_lines[395]		= {inst_bytes[681][0], inst_bytes[681][1], inst_bytes[682][0], inst_bytes[682][1], inst_bytes[682][2], inst_bytes[683][0], inst_bytes[683][1], inst_bytes[683][2]};

		cache_lines[396]		= {inst_bytes[683][3], inst_bytes[683][4], inst_bytes[683][5], inst_bytes[684][0], inst_bytes[684][1], inst_bytes[684][2], inst_bytes[685][0], inst_bytes[685][1]};

		cache_lines[397]		= {inst_bytes[685][2], inst_bytes[685][3], inst_bytes[686][0], inst_bytes[686][1], inst_bytes[686][2], inst_bytes[686][3], inst_bytes[686][4], inst_bytes[686][5]};

		cache_lines[398]		= {inst_bytes[687][0], inst_bytes[687][1], inst_bytes[687][2], inst_bytes[687][3], inst_bytes[687][4], inst_bytes[687][5], inst_bytes[687][6], inst_bytes[688][0]};

		cache_lines[399]		= {inst_bytes[688][1], inst_bytes[689][0], inst_bytes[689][1], inst_bytes[690][0], inst_bytes[690][1], inst_bytes[690][2], inst_bytes[691][0], inst_bytes[691][1]};

		cache_lines[400]		= {inst_bytes[691][2], inst_bytes[691][3], inst_bytes[691][4], inst_bytes[691][5], inst_bytes[692][0], inst_bytes[692][1], inst_bytes[692][2], inst_bytes[693][0]};

		cache_lines[401]		= {inst_bytes[693][1], inst_bytes[693][2], inst_bytes[693][3], inst_bytes[694][0], inst_bytes[694][1], inst_bytes[694][2], inst_bytes[694][3], inst_bytes[694][4]};

		cache_lines[402]		= {inst_bytes[694][5], inst_bytes[695][0], inst_bytes[695][1], inst_bytes[695][2], inst_bytes[695][3], inst_bytes[695][4], inst_bytes[695][5], inst_bytes[695][6]};

		cache_lines[403]		= {inst_bytes[696][0], inst_bytes[696][1], inst_bytes[697][0], inst_bytes[697][1], inst_bytes[697][2], inst_bytes[698][0], inst_bytes[698][1], inst_bytes[698][2]};

		cache_lines[404]		= {inst_bytes[698][3], inst_bytes[699][0], inst_bytes[699][1], inst_bytes[699][2], inst_bytes[699][3], inst_bytes[699][4], inst_bytes[699][5], inst_bytes[699][6]};

		cache_lines[405]		= {inst_bytes[700][0], inst_bytes[700][1], inst_bytes[700][2], inst_bytes[700][3], inst_bytes[701][0], inst_bytes[701][1], inst_bytes[701][2], inst_bytes[701][3]};

		cache_lines[406]		= {inst_bytes[701][4], inst_bytes[702][0], inst_bytes[702][1], inst_bytes[702][2], inst_bytes[702][3], inst_bytes[702][4], inst_bytes[702][5], inst_bytes[702][6]};

		cache_lines[407]		= {inst_bytes[703][0], inst_bytes[703][1], inst_bytes[703][2], inst_bytes[703][3], inst_bytes[703][4], inst_bytes[703][5], inst_bytes[703][6], inst_bytes[703][7]};

		cache_lines[408]		= {inst_bytes[704][0], inst_bytes[704][1], inst_bytes[704][2], inst_bytes[705][0], inst_bytes[705][1], inst_bytes[706][0], inst_bytes[706][1], inst_bytes[706][2]};

		cache_lines[409]		= {inst_bytes[707][0], inst_bytes[707][1], inst_bytes[707][2], inst_bytes[707][3], inst_bytes[707][4], inst_bytes[707][5], inst_bytes[708][0], inst_bytes[708][1]};

		cache_lines[410]		= {inst_bytes[708][2], inst_bytes[709][0], inst_bytes[709][1], inst_bytes[709][2], inst_bytes[709][3], inst_bytes[710][0], inst_bytes[710][1], inst_bytes[710][2]};

		cache_lines[411]		= {inst_bytes[710][3], inst_bytes[710][4], inst_bytes[710][5], inst_bytes[711][0], inst_bytes[711][1], inst_bytes[711][2], inst_bytes[711][3], inst_bytes[711][4]};

		cache_lines[412]		= {inst_bytes[711][5], inst_bytes[711][6], inst_bytes[712][0], inst_bytes[712][1], inst_bytes[713][0], inst_bytes[713][1], inst_bytes[714][0], inst_bytes[714][1]};

		cache_lines[413]		= {inst_bytes[714][2], inst_bytes[715][0], inst_bytes[715][1], inst_bytes[715][2], inst_bytes[715][3], inst_bytes[715][4], inst_bytes[715][5], inst_bytes[716][0]};

		cache_lines[414]		= {inst_bytes[716][1], inst_bytes[716][2], inst_bytes[717][0], inst_bytes[717][1], inst_bytes[717][2], inst_bytes[717][3], inst_bytes[718][0], inst_bytes[718][1]};

		cache_lines[415]		= {inst_bytes[718][2], inst_bytes[718][3], inst_bytes[718][4], inst_bytes[718][5], inst_bytes[719][0], inst_bytes[719][1], inst_bytes[719][2], inst_bytes[719][3]};

		cache_lines[416]		= {inst_bytes[719][4], inst_bytes[719][5], inst_bytes[719][6], inst_bytes[720][0], inst_bytes[720][1], inst_bytes[721][0], inst_bytes[721][1], inst_bytes[721][2]};

		cache_lines[417]		= {inst_bytes[722][0], inst_bytes[722][1], inst_bytes[722][2], inst_bytes[722][3], inst_bytes[723][0], inst_bytes[723][1], inst_bytes[723][2], inst_bytes[723][3]};

		cache_lines[418]		= {inst_bytes[723][4], inst_bytes[723][5], inst_bytes[723][6], inst_bytes[724][0], inst_bytes[724][1], inst_bytes[724][2], inst_bytes[724][3], inst_bytes[725][0]};

		cache_lines[419]		= {inst_bytes[725][1], inst_bytes[725][2], inst_bytes[725][3], inst_bytes[725][4], inst_bytes[726][0], inst_bytes[726][1], inst_bytes[726][2], inst_bytes[726][3]};

		cache_lines[420]		= {inst_bytes[726][4], inst_bytes[726][5], inst_bytes[726][6], inst_bytes[727][0], inst_bytes[727][1], inst_bytes[727][2], inst_bytes[727][3], inst_bytes[727][4]};

		cache_lines[421]		= {inst_bytes[727][5], inst_bytes[727][6], inst_bytes[727][7], inst_bytes[728][0], inst_bytes[728][1], inst_bytes[728][2], inst_bytes[729][0], inst_bytes[729][1]};

		cache_lines[422]		= {inst_bytes[730][0], inst_bytes[730][1], inst_bytes[730][2], inst_bytes[731][0], inst_bytes[731][1], inst_bytes[731][2], inst_bytes[731][3], inst_bytes[731][4]};

		cache_lines[423]		= {inst_bytes[731][5], inst_bytes[732][0], inst_bytes[732][1], inst_bytes[732][2], inst_bytes[733][0], inst_bytes[733][1], inst_bytes[733][2], inst_bytes[733][3]};

		cache_lines[424]		= {inst_bytes[734][0], inst_bytes[734][1], inst_bytes[734][2], inst_bytes[734][3], inst_bytes[734][4], inst_bytes[734][5], inst_bytes[735][0], inst_bytes[735][1]};

		cache_lines[425]		= {inst_bytes[735][2], inst_bytes[735][3], inst_bytes[735][4], inst_bytes[735][5], inst_bytes[735][6], inst_bytes[736][0], inst_bytes[736][1], inst_bytes[737][0]};

		cache_lines[426]		= {inst_bytes[737][1], inst_bytes[738][0], inst_bytes[738][1], inst_bytes[738][2], inst_bytes[739][0], inst_bytes[739][1], inst_bytes[739][2], inst_bytes[739][3]};

		cache_lines[427]		= {inst_bytes[739][4], inst_bytes[739][5], inst_bytes[740][0], inst_bytes[740][1], inst_bytes[740][2], inst_bytes[741][0], inst_bytes[741][1], inst_bytes[741][2]};

		cache_lines[428]		= {inst_bytes[741][3], inst_bytes[742][0], inst_bytes[742][1], inst_bytes[742][2], inst_bytes[742][3], inst_bytes[742][4], inst_bytes[742][5], inst_bytes[743][0]};

		cache_lines[429]		= {inst_bytes[743][1], inst_bytes[743][2], inst_bytes[743][3], inst_bytes[743][4], inst_bytes[743][5], inst_bytes[743][6], inst_bytes[744][0], inst_bytes[744][1]};

		cache_lines[430]		= {inst_bytes[745][0], inst_bytes[745][1], inst_bytes[745][2], inst_bytes[746][0], inst_bytes[746][1], inst_bytes[746][2], inst_bytes[746][3], inst_bytes[747][0]};

		cache_lines[431]		= {inst_bytes[747][1], inst_bytes[747][2], inst_bytes[747][3], inst_bytes[747][4], inst_bytes[747][5], inst_bytes[747][6], inst_bytes[748][0], inst_bytes[748][1]};

		cache_lines[432]		= {inst_bytes[748][2], inst_bytes[748][3], inst_bytes[749][0], inst_bytes[749][1], inst_bytes[749][2], inst_bytes[749][3], inst_bytes[749][4], inst_bytes[750][0]};

		cache_lines[433]		= {inst_bytes[750][1], inst_bytes[750][2], inst_bytes[750][3], inst_bytes[750][4], inst_bytes[750][5], inst_bytes[750][6], inst_bytes[751][0], inst_bytes[751][1]};

		cache_lines[434]		= {inst_bytes[751][2], inst_bytes[751][3], inst_bytes[751][4], inst_bytes[751][5], inst_bytes[751][6], inst_bytes[751][7], inst_bytes[752][0], inst_bytes[752][1]};

		cache_lines[435]		= {inst_bytes[752][2], inst_bytes[753][0], inst_bytes[754][0], inst_bytes[754][1], inst_bytes[755][0], inst_bytes[756][0], inst_bytes[756][1], inst_bytes[757][0]};

		cache_lines[436]		= {inst_bytes[757][1], inst_bytes[757][2], inst_bytes[758][0], inst_bytes[758][1], inst_bytes[758][2], inst_bytes[758][3], inst_bytes[758][4], inst_bytes[758][5]};

		cache_lines[437]		= {inst_bytes[759][0], inst_bytes[759][1], inst_bytes[759][2], inst_bytes[760][0], inst_bytes[760][1], inst_bytes[760][2], inst_bytes[760][3], inst_bytes[761][0]};

		cache_lines[438]		= {inst_bytes[761][1], inst_bytes[761][2], inst_bytes[761][3], inst_bytes[761][4], inst_bytes[761][5], inst_bytes[762][0], inst_bytes[762][1], inst_bytes[762][2]};

		cache_lines[439]		= {inst_bytes[762][3], inst_bytes[762][4], inst_bytes[762][5], inst_bytes[762][6], inst_bytes[763][0], inst_bytes[763][1], inst_bytes[764][0], inst_bytes[764][1]};

		cache_lines[440]		= {inst_bytes[765][0], inst_bytes[765][1], inst_bytes[765][2], inst_bytes[766][0], inst_bytes[766][1], inst_bytes[766][2], inst_bytes[766][3], inst_bytes[766][4]};

		cache_lines[441]		= {inst_bytes[766][5], inst_bytes[767][0], inst_bytes[767][1], inst_bytes[767][2], inst_bytes[768][0], inst_bytes[768][1], inst_bytes[768][2], inst_bytes[768][3]};

		cache_lines[442]		= {inst_bytes[769][0], inst_bytes[769][1], inst_bytes[769][2], inst_bytes[769][3], inst_bytes[769][4], inst_bytes[769][5], inst_bytes[770][0], inst_bytes[770][1]};

		cache_lines[443]		= {inst_bytes[770][2], inst_bytes[770][3], inst_bytes[770][4], inst_bytes[770][5], inst_bytes[770][6], inst_bytes[771][0], inst_bytes[771][1], inst_bytes[772][0]};

		cache_lines[444]		= {inst_bytes[772][1], inst_bytes[773][0], inst_bytes[773][1], inst_bytes[773][2], inst_bytes[774][0], inst_bytes[774][1], inst_bytes[774][2], inst_bytes[774][3]};

		cache_lines[445]		= {inst_bytes[774][4], inst_bytes[774][5], inst_bytes[775][0], inst_bytes[775][1], inst_bytes[775][2], inst_bytes[776][0], inst_bytes[776][1], inst_bytes[776][2]};

		cache_lines[446]		= {inst_bytes[776][3], inst_bytes[777][0], inst_bytes[777][1], inst_bytes[777][2], inst_bytes[777][3], inst_bytes[777][4], inst_bytes[777][5], inst_bytes[778][0]};

		cache_lines[447]		= {inst_bytes[778][1], inst_bytes[778][2], inst_bytes[778][3], inst_bytes[778][4], inst_bytes[778][5], inst_bytes[778][6], inst_bytes[779][0], inst_bytes[779][1]};
	end
	//Fetch 
	reg		[0:0]	CLK;
	reg		[0:0]	reset;
	
	reg		[63:0]	cache_line;
	reg		[0:0]	cache_line_valid;
	wire	[43:0]	tlb_trans;
	wire	[0:0]	tlb_hit;
	wire	[31:0]	bpred_target;
	wire	[0:0]	bpred_taken;
	wire	[0:0]	bpred_hit;
	wire	[0:0]	dec1_stall;
	reg		[0:0]	data_gp_excp;
	reg		[0:0]	data_pf_excp;
	reg		[31:0]	data_excp_eip;
	reg		[31:0]	ex_branch_eip;
	reg		[31:0]	ex_branch_target;
	reg		[0:0]	ex_branch_taken;
	reg		[0:0]	ex_branch_mispred;
	reg		[0:0]	ex_branch_valid;
	reg		[15:0] 	cs_in;
	reg		[0:0] 	cs_en;
	reg		[7:0]	intr_vec;
	
	wire	[0:0]	replay_inst;
	reg		[31:0]	replay_eip;
	
	
	wire	[31:0]	fetch_addr;
	wire	[0:0]	fetch_addr_valid;
	wire	[31:0]	tlb_addr;
	wire	[0:0]	tlb_access;
	wire	[31:0]	bpred_pc_out;
	wire	[31:0]	update_bpred_pc;
	wire	[31:0]	update_bpred_target;
	wire	[0:0]	update_bpred_taken;
	wire	[0:0]	update_bpred_valid;
	wire	[63:0]	fetch_bytes;
	wire	[255:0]	fetch_pcs;
	wire	[0:0]	fetch_not_ready;
	wire	[3:0]	fetch_width;
	wire	[0:0]	page_bound;
	wire	[3:0]	br_fetch_id;
	wire	[31:0]	fetch_bpred_tgt;
	wire	[0:0]	fetch_bpred_taken;
	wire	[0:0]	fetch_ex_br_taken;
	
	//Decode1
	wire	[0:0]	has_prefix1;
	wire	[0:0]	has_prefix2;
	wire	[0:0]	has_prefix3;
	wire	[0:0]	has_op2;
	wire	[0:0]	has_imm8;
	wire	[0:0]	has_imm16;
	wire	[0:0]	has_imm32;
	wire	[0:0]	has_modrm;
	wire	[0:0]	has_sib;
	wire	[0:0]	has_disp8;
	wire	[0:0]	has_disp32;
	wire	[7:0]	prefix2_byte;
	wire	[7:0]	opcode1_byte;
	wire	[7:0]	opcode2_byte;
	wire	[7:0]	modrm_byte;
	wire	[7:0]	sib_byte;
	wire	[3:0]	size;
	wire	[7:0]	b0_out;
	wire	[7:0]	b1_out;
	wire	[7:0]	b2_out;
	wire	[7:0]	b3_out;
	wire	[7:0]	b4_out;
	wire	[7:0]	b5_out;
	wire	[7:0]	b6_out;
	wire	[7:0]	b7_out;
	wire	[7:0]	b8_out;
	wire	[7:0]	b9_out;
	wire	[7:0]	b10_out;
	wire	[7:0]	b11_out;
	wire	[7:0]	b12_out;
	
	wire	[0:0]	dec2_stall;
	wire	[31:0]	eip;
	wire	[31:0]	n_eip;
	wire	[0:0]	dec1_not_ready;
	wire	[3:0]	br_fetch_id_out;
	wire	[31:0]	d1_bpred_tgt;
	wire	[0:0]	d1_bpred_taken;
	wire	[0:0]	d1_ex_br_taken;
	
	
	fetch 			ft(	CLK, 
						reset, 
						cache_line, 
						cache_line_valid,
						tlb_trans,
						tlb_hit,
						bpred_target,
						bpred_taken, 
						bpred_hit,
						dec1_stall,
						replay_inst,
						replay_eip,
						data_gp_excp,
						data_pf_excp,
						data_excp_eip,
						ex_branch_eip,
						ex_branch_target, 
						ex_branch_taken,
						ex_branch_mispred,						
						ex_branch_valid,
						cs_in,
						cs_en,
						intr_vec,
						
						fetch_addr,
						fetch_addr_valid,
						tlb_addr, 
						tlb_access, 
						bpred_pc_out, 
						update_bpred_pc,
						update_bpred_target,
						update_bpred_taken,
						update_bpred_mispred,
						update_bpred_valid,
						fetch_bytes,
						fetch_pcs,
						fetch_not_ready,
						fetch_width,
						page_bound,
						br_fetch_id,
						fetch_bpred_tgt,
						fetch_bpred_taken,
						fetch_ex_br_taken
						);
						
	reg		[351:0]		tlb_init;
	tlb				mtlb(
						tlb_addr, 
						tlb_access,
						tlb_trans,
						tlb_hit,
						,
						,
						,
						,
						tlb_init);
						
						
	bpred 			br	(
						CLK,
						reset,
						bpred_pc_out,
						
						update_bpred_pc,
						update_bpred_target,
						update_bpred_taken,
						update_bpred_mispred,
						update_bpred_valid,
						
						bpred_target,
						bpred_taken,
						bpred_hit
						);
	
	wire	[0:0]	bytes_cleanup;
	wire	[3:0]	cleanup_id;	
	reg		[0:0]	datapath_inv;
	
	decode1			d1(	CLK, 
						reset, 
						{fetch_ex_br_taken, fetch_bpred_taken, fetch_bpred_tgt, br_fetch_id, fetch_pcs[31:0], fetch_bytes[7:0]},
						{fetch_ex_br_taken, fetch_bpred_taken, fetch_bpred_tgt, br_fetch_id, fetch_pcs[63:32], fetch_bytes[15:8]},
						{fetch_ex_br_taken, fetch_bpred_taken, fetch_bpred_tgt, br_fetch_id, fetch_pcs[95:64], fetch_bytes[23:16]},
						{fetch_ex_br_taken, fetch_bpred_taken, fetch_bpred_tgt, br_fetch_id, fetch_pcs[127:96], fetch_bytes[31:24]},
						{fetch_ex_br_taken, fetch_bpred_taken, fetch_bpred_tgt, br_fetch_id, fetch_pcs[159:128], fetch_bytes[39:32]},
						{fetch_ex_br_taken, fetch_bpred_taken, fetch_bpred_tgt, br_fetch_id, fetch_pcs[191:160], fetch_bytes[47:40]},
						{fetch_ex_br_taken, fetch_bpred_taken, fetch_bpred_tgt, br_fetch_id, fetch_pcs[223:192], fetch_bytes[55:48]},
						{fetch_ex_br_taken, fetch_bpred_taken, fetch_bpred_tgt, br_fetch_id, fetch_pcs[255:224], fetch_bytes[63:56]},
						dec2_stall, 
						fetch_not_ready,
						fetch_width,
						page_bound,
						bytes_cleanup,
						cleanup_id,
						datapath_inv, 
						replay_inst,
						
						has_prefix1, 
						has_prefix2, 
						has_prefix3, 
						has_op2, 
						has_imm8, 
						has_imm16, 
						has_imm32, 
						has_modrm, 
						has_sib, 
						has_disp8, 
						has_disp32, 
						size,
						prefix2_byte, 
						opcode1_byte, 
						opcode2_byte, 
						modrm_byte, 
						sib_byte, 
						b0_out, 
						b1_out, 
						b2_out, 
						b3_out, 
						b4_out, 
						b5_out, 
						b6_out, 
						b7_out, 
						b8_out, 
						b9_out, 
						b10_out, 
						b11_out, 
						b12_out, 
						eip,
						dec1_stall, 
						dec1_not_ready,
						br_fetch_id_out,
						d1_bpred_tgt,
						d1_bpred_taken,
						d1_ex_br_taken
						);
	
	reg [0:0]  rr_stall; 
	wire [59:0] i_CS;        
	wire [31:0] i_imm;       
	wire [31:0] i_disp;
	wire [1:0] i_immSize;       
	wire [1:0] i_dispSize;	
	wire [0:0]	i_SIB;
	wire [1:0]  i_scale;    
	wire [0:0]  i_baseRen;      
	wire [0:0]  i_idxRen;        
	wire [31:0] i_nEIP;      
	wire [31:0] i_EIP;       
	wire [31:0] i_bp_tgt;    
	wire [15:0] i_currCS;    
	wire [7:0]  i_imm8;      
	wire [1:0]  i_opSize;   
	wire [2:0]  i_sr1;       
	wire [2:0]  i_sr2;       
	wire [2:0]  i_base;      
	wire [2:0]  i_idx;       
	wire [2:0]  i_segR1;     
	wire [2:0]  i_segR2;     
	wire [0:0]  i_bp_taken;  
	wire [0:0]  i_indir_addr;     
	wire [0:0]  i_Dflag;     
	wire [0:0]  i_v;
	wire [3:0]  i_br_fetch_id;
						
	decode2			d2(	CLK,
						reset,
						
						has_prefix1,
						has_prefix2,
						has_prefix3,
						has_imm8,
						has_imm16,
						has_imm32,
						has_disp8,
						has_disp32,
						has_op2,
						has_modrm,
						has_sib,
						
						size,
						
						prefix2_byte,
						opcode1_byte,
						opcode2_byte,
						modrm_byte,
						sib_byte,
						
						b0_out,
						b1_out,
						b2_out,
						b3_out,
						b4_out,
						b5_out,
						b6_out,
						b7_out,
						b8_out,
						b9_out,
						b10_out,
						b11_out,
						b12_out,
						
						eip,
						dec1_not_ready,
						br_fetch_id_out,
						d1_bpred_tgt,
						d1_bpred_taken,
						d1_ex_br_taken,
						
						rr_stall,
						
						dec2_stall,
						bytes_cleanup,
						cleanup_id,
						replay_inst,
						
						//Pipeline read reg
						i_CS,			i_imm,		i_disp,      
						i_immSize,		i_dispSize, i_SIB,
						i_scale,		i_baseRen, 	i_idxRen,
						i_nEIP,			i_EIP,		i_bp_tgt,    
						i_imm8,			i_opSize,	i_sr1,
						i_sr2,			i_base,		i_idx,
						i_segR1,		i_segR2,	i_bp_taken,
						i_indir_addr,	i_Dflag,    i_br_fetch_id, 
						i_v 		  
						);
						
	
	always
	begin
		#6 CLK = !CLK;
	end
	
	
	//Assertions
	integer i = 0;
	always@ (posedge CLK)
	begin
	
		
		if(!dec1_not_ready && !dec2_stall)
		begin
			if(inst_size[i]!=size) 
			begin
				$display("Error. Index=%d, calc_size=%d, actual_size=%d\n", i, size, inst_size[i]);
			end
			i = i + 1;
			if(i==780)
			begin
				i = 0;
				$fclose(f);
				$finish;
			end
		end
	
	end

	integer f;
	always@ (posedge CLK)
	begin
		if(i_v)
		begin
			$fwrite(f, "%b\n", i_CS);
		end
	end

	initial begin
	
		f = $fopen("control_out", "w");
		CLK = 0;
		reset = 0;
		
		$readmemb("cs_bits.mem", d2.cs.rm.rm0h.mem);
		$readmemb("./cs_files/cs0_l.mem", d2.cs.rm.rm0l.mem);
		$readmemb("cs_bits.mem", d2.cs.rm.rm1h.mem);
		$readmemb("./cs_files/cs1_l.mem", d2.cs.rm.rm1l.mem);
		$readmemb("cs_bits.mem", d2.cs.rm.rm2h.mem);
		$readmemb("./cs_files/cs2_l.mem", d2.cs.rm.rm2l.mem);
		$readmemb("cs_bits.mem", d2.cs.rm.rm3h.mem);
		$readmemb("./cs_files/cs3_l.mem", d2.cs.rm.rm3l.mem);
		$readmemb("cs_bits.mem", d2.cs.rm.rm4h.mem);
		$readmemb("./cs_files/cs4_l.mem", d2.cs.rm.rm4l.mem);
		$readmemb("cs_bits.mem", d2.cs.rm.rm5h.mem);
		$readmemb("./cs_files/cs5_l.mem", d2.cs.rm.rm5l.mem);
		$readmemb("cs_bits.mem", d2.cs.rm.rm6h.mem);
		$readmemb("./cs_files/cs6_l.mem", d2.cs.rm.rm6l.mem);
		$readmemb("cs_bits.mem", d2.cs.rm.rm7h.mem);
		$readmemb("./cs_files/cs7_l.mem", d2.cs.rm.rm7l.mem);
		
		
		cache_line 			= 63'h0;
		cache_line_valid 	= 0;
		
		data_gp_excp 		= 1'b0;
		data_pf_excp 		= 1'b0;
		data_excp_eip		= 32'b0;
		ex_branch_eip 		= 32'b0;
		ex_branch_target	= 32'b0;
		ex_branch_taken		= 1'b0;
		ex_branch_mispred	= 1'b0;
		ex_branch_valid		= 1'b0;
		intr_vec			= 8'b0;
		datapath_inv		= 1'b0;
		
		cs_in				= 1'b0;
		cs_en				= 1'b0;
		
		replay_eip			= 32'd0;
		rr_stall			= 1'b0;
		tlb_init			= {{1'b1, 20'h0,20'h1,1'b1,1'b1,1'b0}, {1'b1, 20'h2000,20'h2,1'b1,1'b1,1'b1}, {1'b1, 20'h4000,20'h5,1'b1,1'b1,1'b1}, {1'b1, 20'hb000,20'h4,1'b1,1'b1,1'b1}, {1'b1, 20'hc000,20'h7,1'b1,1'b1,1'b1}, {1'b1, 20'ha000,20'h5,1'b1,1'b1,1'b1}, {1'b1, 20'h8000,20'h1,1'b1,1'b1,1'b1}, {1'b1, 20'h9000,20'h3,1'b1,1'b1,1'b1}};
	
		#13.5
		reset 				= 1;
		cache_line_valid	= 1'b0;


	end
	
	integer j = 0;
	//Feed cache lines
	always@(reset, fetch_addr_valid, fetch_addr)
	begin
		if(reset==1'b1 && fetch_addr_valid==1'b1)
		begin
			cache_line_valid	= 1'b1;
			cache_line = cache_lines[(fetch_addr[11:0]>>3)];
			//if(j==448)
			//begin
				//cache_line_valid = 1'b0;
			//	j = 0;
			//end
		end
	end
	
	
endmodule